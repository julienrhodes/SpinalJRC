-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2017.08.27940

-- Build Date:         Sep 12 2017 08:26:01

-- File Generated:     Apr 28 2020 10:13:15

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "MyTopLevel" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of MyTopLevel
entity MyTopLevel is
port (
    io_leds : out std_logic_vector(7 downto 0);
    io_jtag_tms : in std_logic;
    io_jtag_tdo : out std_logic;
    io_jtag_tdi : in std_logic;
    io_jtag_tck : in std_logic;
    global_reset : in std_logic;
    global_clk : in std_logic);
end MyTopLevel;

-- Architecture of MyTopLevel
-- View name is \INTERFACE\
architecture \INTERFACE\ of MyTopLevel is

signal \N__5400\ : std_logic;
signal \N__5399\ : std_logic;
signal \N__5398\ : std_logic;
signal \N__5389\ : std_logic;
signal \N__5388\ : std_logic;
signal \N__5387\ : std_logic;
signal \N__5380\ : std_logic;
signal \N__5379\ : std_logic;
signal \N__5378\ : std_logic;
signal \N__5371\ : std_logic;
signal \N__5370\ : std_logic;
signal \N__5369\ : std_logic;
signal \N__5362\ : std_logic;
signal \N__5361\ : std_logic;
signal \N__5360\ : std_logic;
signal \N__5353\ : std_logic;
signal \N__5352\ : std_logic;
signal \N__5351\ : std_logic;
signal \N__5344\ : std_logic;
signal \N__5343\ : std_logic;
signal \N__5342\ : std_logic;
signal \N__5335\ : std_logic;
signal \N__5334\ : std_logic;
signal \N__5333\ : std_logic;
signal \N__5326\ : std_logic;
signal \N__5325\ : std_logic;
signal \N__5324\ : std_logic;
signal \N__5317\ : std_logic;
signal \N__5316\ : std_logic;
signal \N__5315\ : std_logic;
signal \N__5308\ : std_logic;
signal \N__5307\ : std_logic;
signal \N__5306\ : std_logic;
signal \N__5299\ : std_logic;
signal \N__5298\ : std_logic;
signal \N__5297\ : std_logic;
signal \N__5290\ : std_logic;
signal \N__5289\ : std_logic;
signal \N__5288\ : std_logic;
signal \N__5281\ : std_logic;
signal \N__5280\ : std_logic;
signal \N__5279\ : std_logic;
signal \N__5262\ : std_logic;
signal \N__5261\ : std_logic;
signal \N__5258\ : std_logic;
signal \N__5257\ : std_logic;
signal \N__5254\ : std_logic;
signal \N__5251\ : std_logic;
signal \N__5248\ : std_logic;
signal \N__5245\ : std_logic;
signal \N__5238\ : std_logic;
signal \N__5235\ : std_logic;
signal \N__5232\ : std_logic;
signal \N__5229\ : std_logic;
signal \N__5228\ : std_logic;
signal \N__5225\ : std_logic;
signal \N__5222\ : std_logic;
signal \N__5217\ : std_logic;
signal \N__5216\ : std_logic;
signal \N__5215\ : std_logic;
signal \N__5214\ : std_logic;
signal \N__5213\ : std_logic;
signal \N__5202\ : std_logic;
signal \N__5199\ : std_logic;
signal \N__5196\ : std_logic;
signal \N__5195\ : std_logic;
signal \N__5192\ : std_logic;
signal \N__5189\ : std_logic;
signal \N__5186\ : std_logic;
signal \N__5185\ : std_logic;
signal \N__5182\ : std_logic;
signal \N__5181\ : std_logic;
signal \N__5178\ : std_logic;
signal \N__5175\ : std_logic;
signal \N__5172\ : std_logic;
signal \N__5169\ : std_logic;
signal \N__5164\ : std_logic;
signal \N__5157\ : std_logic;
signal \N__5154\ : std_logic;
signal \N__5151\ : std_logic;
signal \N__5148\ : std_logic;
signal \N__5145\ : std_logic;
signal \N__5144\ : std_logic;
signal \N__5141\ : std_logic;
signal \N__5138\ : std_logic;
signal \N__5133\ : std_logic;
signal \N__5132\ : std_logic;
signal \N__5127\ : std_logic;
signal \N__5124\ : std_logic;
signal \N__5121\ : std_logic;
signal \N__5120\ : std_logic;
signal \N__5115\ : std_logic;
signal \N__5112\ : std_logic;
signal \N__5109\ : std_logic;
signal \N__5106\ : std_logic;
signal \N__5103\ : std_logic;
signal \N__5102\ : std_logic;
signal \N__5099\ : std_logic;
signal \N__5096\ : std_logic;
signal \N__5091\ : std_logic;
signal \N__5090\ : std_logic;
signal \N__5085\ : std_logic;
signal \N__5082\ : std_logic;
signal \N__5079\ : std_logic;
signal \N__5078\ : std_logic;
signal \N__5077\ : std_logic;
signal \N__5076\ : std_logic;
signal \N__5075\ : std_logic;
signal \N__5074\ : std_logic;
signal \N__5071\ : std_logic;
signal \N__5068\ : std_logic;
signal \N__5065\ : std_logic;
signal \N__5064\ : std_logic;
signal \N__5063\ : std_logic;
signal \N__5062\ : std_logic;
signal \N__5061\ : std_logic;
signal \N__5058\ : std_logic;
signal \N__5057\ : std_logic;
signal \N__5056\ : std_logic;
signal \N__5055\ : std_logic;
signal \N__5054\ : std_logic;
signal \N__5053\ : std_logic;
signal \N__5052\ : std_logic;
signal \N__5051\ : std_logic;
signal \N__5050\ : std_logic;
signal \N__5049\ : std_logic;
signal \N__5048\ : std_logic;
signal \N__5047\ : std_logic;
signal \N__5046\ : std_logic;
signal \N__5045\ : std_logic;
signal \N__5044\ : std_logic;
signal \N__5043\ : std_logic;
signal \N__5042\ : std_logic;
signal \N__5041\ : std_logic;
signal \N__5040\ : std_logic;
signal \N__5039\ : std_logic;
signal \N__5038\ : std_logic;
signal \N__5037\ : std_logic;
signal \N__5032\ : std_logic;
signal \N__5027\ : std_logic;
signal \N__5024\ : std_logic;
signal \N__5021\ : std_logic;
signal \N__5014\ : std_logic;
signal \N__5011\ : std_logic;
signal \N__5002\ : std_logic;
signal \N__4991\ : std_logic;
signal \N__4986\ : std_logic;
signal \N__4979\ : std_logic;
signal \N__4968\ : std_logic;
signal \N__4963\ : std_logic;
signal \N__4956\ : std_logic;
signal \N__4951\ : std_logic;
signal \N__4944\ : std_logic;
signal \N__4929\ : std_logic;
signal \N__4928\ : std_logic;
signal \N__4927\ : std_logic;
signal \N__4926\ : std_logic;
signal \N__4925\ : std_logic;
signal \N__4924\ : std_logic;
signal \N__4923\ : std_logic;
signal \N__4922\ : std_logic;
signal \N__4921\ : std_logic;
signal \N__4920\ : std_logic;
signal \N__4919\ : std_logic;
signal \N__4918\ : std_logic;
signal \N__4917\ : std_logic;
signal \N__4916\ : std_logic;
signal \N__4915\ : std_logic;
signal \N__4914\ : std_logic;
signal \N__4913\ : std_logic;
signal \N__4912\ : std_logic;
signal \N__4911\ : std_logic;
signal \N__4910\ : std_logic;
signal \N__4907\ : std_logic;
signal \N__4906\ : std_logic;
signal \N__4905\ : std_logic;
signal \N__4904\ : std_logic;
signal \N__4901\ : std_logic;
signal \N__4900\ : std_logic;
signal \N__4899\ : std_logic;
signal \N__4898\ : std_logic;
signal \N__4897\ : std_logic;
signal \N__4896\ : std_logic;
signal \N__4885\ : std_logic;
signal \N__4878\ : std_logic;
signal \N__4877\ : std_logic;
signal \N__4874\ : std_logic;
signal \N__4871\ : std_logic;
signal \N__4870\ : std_logic;
signal \N__4867\ : std_logic;
signal \N__4866\ : std_logic;
signal \N__4865\ : std_logic;
signal \N__4864\ : std_logic;
signal \N__4863\ : std_logic;
signal \N__4860\ : std_logic;
signal \N__4859\ : std_logic;
signal \N__4858\ : std_logic;
signal \N__4857\ : std_logic;
signal \N__4856\ : std_logic;
signal \N__4855\ : std_logic;
signal \N__4854\ : std_logic;
signal \N__4851\ : std_logic;
signal \N__4848\ : std_logic;
signal \N__4841\ : std_logic;
signal \N__4832\ : std_logic;
signal \N__4825\ : std_logic;
signal \N__4822\ : std_logic;
signal \N__4815\ : std_logic;
signal \N__4810\ : std_logic;
signal \N__4807\ : std_logic;
signal \N__4804\ : std_logic;
signal \N__4801\ : std_logic;
signal \N__4796\ : std_logic;
signal \N__4791\ : std_logic;
signal \N__4786\ : std_logic;
signal \N__4779\ : std_logic;
signal \N__4770\ : std_logic;
signal \N__4767\ : std_logic;
signal \N__4758\ : std_logic;
signal \N__4751\ : std_logic;
signal \N__4728\ : std_logic;
signal \N__4727\ : std_logic;
signal \N__4724\ : std_logic;
signal \N__4719\ : std_logic;
signal \N__4716\ : std_logic;
signal \N__4715\ : std_logic;
signal \N__4714\ : std_logic;
signal \N__4713\ : std_logic;
signal \N__4712\ : std_logic;
signal \N__4711\ : std_logic;
signal \N__4710\ : std_logic;
signal \N__4709\ : std_logic;
signal \N__4708\ : std_logic;
signal \N__4707\ : std_logic;
signal \N__4706\ : std_logic;
signal \N__4705\ : std_logic;
signal \N__4704\ : std_logic;
signal \N__4703\ : std_logic;
signal \N__4702\ : std_logic;
signal \N__4701\ : std_logic;
signal \N__4700\ : std_logic;
signal \N__4665\ : std_logic;
signal \N__4662\ : std_logic;
signal \N__4659\ : std_logic;
signal \N__4656\ : std_logic;
signal \N__4653\ : std_logic;
signal \N__4650\ : std_logic;
signal \N__4649\ : std_logic;
signal \N__4646\ : std_logic;
signal \N__4643\ : std_logic;
signal \N__4640\ : std_logic;
signal \N__4637\ : std_logic;
signal \N__4636\ : std_logic;
signal \N__4631\ : std_logic;
signal \N__4628\ : std_logic;
signal \N__4623\ : std_logic;
signal \N__4622\ : std_logic;
signal \N__4619\ : std_logic;
signal \N__4616\ : std_logic;
signal \N__4613\ : std_logic;
signal \N__4610\ : std_logic;
signal \N__4605\ : std_logic;
signal \N__4602\ : std_logic;
signal \N__4599\ : std_logic;
signal \N__4596\ : std_logic;
signal \N__4595\ : std_logic;
signal \N__4592\ : std_logic;
signal \N__4589\ : std_logic;
signal \N__4588\ : std_logic;
signal \N__4583\ : std_logic;
signal \N__4580\ : std_logic;
signal \N__4575\ : std_logic;
signal \N__4572\ : std_logic;
signal \N__4571\ : std_logic;
signal \N__4568\ : std_logic;
signal \N__4565\ : std_logic;
signal \N__4560\ : std_logic;
signal \N__4557\ : std_logic;
signal \N__4554\ : std_logic;
signal \N__4551\ : std_logic;
signal \N__4548\ : std_logic;
signal \N__4545\ : std_logic;
signal \N__4544\ : std_logic;
signal \N__4541\ : std_logic;
signal \N__4538\ : std_logic;
signal \N__4537\ : std_logic;
signal \N__4532\ : std_logic;
signal \N__4529\ : std_logic;
signal \N__4524\ : std_logic;
signal \N__4521\ : std_logic;
signal \N__4520\ : std_logic;
signal \N__4517\ : std_logic;
signal \N__4514\ : std_logic;
signal \N__4511\ : std_logic;
signal \N__4508\ : std_logic;
signal \N__4503\ : std_logic;
signal \N__4500\ : std_logic;
signal \N__4497\ : std_logic;
signal \N__4496\ : std_logic;
signal \N__4493\ : std_logic;
signal \N__4490\ : std_logic;
signal \N__4485\ : std_logic;
signal \N__4482\ : std_logic;
signal \N__4481\ : std_logic;
signal \N__4478\ : std_logic;
signal \N__4475\ : std_logic;
signal \N__4472\ : std_logic;
signal \N__4469\ : std_logic;
signal \N__4464\ : std_logic;
signal \N__4461\ : std_logic;
signal \N__4458\ : std_logic;
signal \N__4457\ : std_logic;
signal \N__4454\ : std_logic;
signal \N__4451\ : std_logic;
signal \N__4450\ : std_logic;
signal \N__4447\ : std_logic;
signal \N__4444\ : std_logic;
signal \N__4441\ : std_logic;
signal \N__4434\ : std_logic;
signal \N__4431\ : std_logic;
signal \N__4428\ : std_logic;
signal \N__4427\ : std_logic;
signal \N__4424\ : std_logic;
signal \N__4421\ : std_logic;
signal \N__4416\ : std_logic;
signal \N__4413\ : std_logic;
signal \N__4412\ : std_logic;
signal \N__4409\ : std_logic;
signal \N__4408\ : std_logic;
signal \N__4405\ : std_logic;
signal \N__4402\ : std_logic;
signal \N__4399\ : std_logic;
signal \N__4392\ : std_logic;
signal \N__4389\ : std_logic;
signal \N__4388\ : std_logic;
signal \N__4385\ : std_logic;
signal \N__4382\ : std_logic;
signal \N__4379\ : std_logic;
signal \N__4376\ : std_logic;
signal \N__4371\ : std_logic;
signal \N__4368\ : std_logic;
signal \N__4367\ : std_logic;
signal \N__4366\ : std_logic;
signal \N__4365\ : std_logic;
signal \N__4364\ : std_logic;
signal \N__4363\ : std_logic;
signal \N__4362\ : std_logic;
signal \N__4361\ : std_logic;
signal \N__4358\ : std_logic;
signal \N__4343\ : std_logic;
signal \N__4342\ : std_logic;
signal \N__4341\ : std_logic;
signal \N__4338\ : std_logic;
signal \N__4335\ : std_logic;
signal \N__4330\ : std_logic;
signal \N__4323\ : std_logic;
signal \N__4320\ : std_logic;
signal \N__4317\ : std_logic;
signal \N__4314\ : std_logic;
signal \N__4313\ : std_logic;
signal \N__4310\ : std_logic;
signal \N__4307\ : std_logic;
signal \N__4306\ : std_logic;
signal \N__4303\ : std_logic;
signal \N__4300\ : std_logic;
signal \N__4297\ : std_logic;
signal \N__4290\ : std_logic;
signal \N__4289\ : std_logic;
signal \N__4288\ : std_logic;
signal \N__4287\ : std_logic;
signal \N__4286\ : std_logic;
signal \N__4285\ : std_logic;
signal \N__4284\ : std_logic;
signal \N__4283\ : std_logic;
signal \N__4274\ : std_logic;
signal \N__4265\ : std_logic;
signal \N__4260\ : std_logic;
signal \N__4257\ : std_logic;
signal \N__4254\ : std_logic;
signal \N__4253\ : std_logic;
signal \N__4250\ : std_logic;
signal \N__4247\ : std_logic;
signal \N__4244\ : std_logic;
signal \N__4241\ : std_logic;
signal \N__4236\ : std_logic;
signal \N__4233\ : std_logic;
signal \N__4230\ : std_logic;
signal \N__4227\ : std_logic;
signal \N__4224\ : std_logic;
signal \N__4223\ : std_logic;
signal \N__4222\ : std_logic;
signal \N__4221\ : std_logic;
signal \N__4220\ : std_logic;
signal \N__4219\ : std_logic;
signal \N__4218\ : std_logic;
signal \N__4217\ : std_logic;
signal \N__4216\ : std_logic;
signal \N__4215\ : std_logic;
signal \N__4214\ : std_logic;
signal \N__4213\ : std_logic;
signal \N__4210\ : std_logic;
signal \N__4195\ : std_logic;
signal \N__4192\ : std_logic;
signal \N__4189\ : std_logic;
signal \N__4188\ : std_logic;
signal \N__4185\ : std_logic;
signal \N__4184\ : std_logic;
signal \N__4183\ : std_logic;
signal \N__4182\ : std_logic;
signal \N__4179\ : std_logic;
signal \N__4178\ : std_logic;
signal \N__4177\ : std_logic;
signal \N__4176\ : std_logic;
signal \N__4175\ : std_logic;
signal \N__4174\ : std_logic;
signal \N__4173\ : std_logic;
signal \N__4172\ : std_logic;
signal \N__4171\ : std_logic;
signal \N__4170\ : std_logic;
signal \N__4169\ : std_logic;
signal \N__4168\ : std_logic;
signal \N__4161\ : std_logic;
signal \N__4158\ : std_logic;
signal \N__4151\ : std_logic;
signal \N__4148\ : std_logic;
signal \N__4147\ : std_logic;
signal \N__4146\ : std_logic;
signal \N__4141\ : std_logic;
signal \N__4138\ : std_logic;
signal \N__4127\ : std_logic;
signal \N__4116\ : std_logic;
signal \N__4111\ : std_logic;
signal \N__4106\ : std_logic;
signal \N__4101\ : std_logic;
signal \N__4086\ : std_logic;
signal \N__4085\ : std_logic;
signal \N__4084\ : std_logic;
signal \N__4083\ : std_logic;
signal \N__4080\ : std_logic;
signal \N__4077\ : std_logic;
signal \N__4076\ : std_logic;
signal \N__4073\ : std_logic;
signal \N__4072\ : std_logic;
signal \N__4071\ : std_logic;
signal \N__4070\ : std_logic;
signal \N__4069\ : std_logic;
signal \N__4068\ : std_logic;
signal \N__4067\ : std_logic;
signal \N__4066\ : std_logic;
signal \N__4065\ : std_logic;
signal \N__4064\ : std_logic;
signal \N__4063\ : std_logic;
signal \N__4062\ : std_logic;
signal \N__4059\ : std_logic;
signal \N__4054\ : std_logic;
signal \N__4053\ : std_logic;
signal \N__4052\ : std_logic;
signal \N__4051\ : std_logic;
signal \N__4048\ : std_logic;
signal \N__4045\ : std_logic;
signal \N__4042\ : std_logic;
signal \N__4039\ : std_logic;
signal \N__4038\ : std_logic;
signal \N__4033\ : std_logic;
signal \N__4030\ : std_logic;
signal \N__4023\ : std_logic;
signal \N__4014\ : std_logic;
signal \N__4011\ : std_logic;
signal \N__4004\ : std_logic;
signal \N__3997\ : std_logic;
signal \N__3992\ : std_logic;
signal \N__3975\ : std_logic;
signal \N__3974\ : std_logic;
signal \N__3973\ : std_logic;
signal \N__3972\ : std_logic;
signal \N__3969\ : std_logic;
signal \N__3968\ : std_logic;
signal \N__3965\ : std_logic;
signal \N__3964\ : std_logic;
signal \N__3963\ : std_logic;
signal \N__3962\ : std_logic;
signal \N__3961\ : std_logic;
signal \N__3958\ : std_logic;
signal \N__3955\ : std_logic;
signal \N__3950\ : std_logic;
signal \N__3945\ : std_logic;
signal \N__3938\ : std_logic;
signal \N__3937\ : std_logic;
signal \N__3934\ : std_logic;
signal \N__3933\ : std_logic;
signal \N__3930\ : std_logic;
signal \N__3923\ : std_logic;
signal \N__3920\ : std_logic;
signal \N__3917\ : std_logic;
signal \N__3914\ : std_logic;
signal \N__3909\ : std_logic;
signal \N__3906\ : std_logic;
signal \N__3903\ : std_logic;
signal \N__3900\ : std_logic;
signal \N__3897\ : std_logic;
signal \N__3894\ : std_logic;
signal \N__3889\ : std_logic;
signal \N__3882\ : std_logic;
signal \N__3881\ : std_logic;
signal \N__3880\ : std_logic;
signal \N__3875\ : std_logic;
signal \N__3872\ : std_logic;
signal \N__3871\ : std_logic;
signal \N__3870\ : std_logic;
signal \N__3869\ : std_logic;
signal \N__3868\ : std_logic;
signal \N__3865\ : std_logic;
signal \N__3864\ : std_logic;
signal \N__3863\ : std_logic;
signal \N__3862\ : std_logic;
signal \N__3861\ : std_logic;
signal \N__3860\ : std_logic;
signal \N__3859\ : std_logic;
signal \N__3858\ : std_logic;
signal \N__3857\ : std_logic;
signal \N__3856\ : std_logic;
signal \N__3855\ : std_logic;
signal \N__3854\ : std_logic;
signal \N__3853\ : std_logic;
signal \N__3850\ : std_logic;
signal \N__3843\ : std_logic;
signal \N__3840\ : std_logic;
signal \N__3839\ : std_logic;
signal \N__3838\ : std_logic;
signal \N__3835\ : std_logic;
signal \N__3832\ : std_logic;
signal \N__3829\ : std_logic;
signal \N__3818\ : std_logic;
signal \N__3807\ : std_logic;
signal \N__3800\ : std_logic;
signal \N__3795\ : std_logic;
signal \N__3780\ : std_logic;
signal \N__3777\ : std_logic;
signal \N__3774\ : std_logic;
signal \N__3771\ : std_logic;
signal \N__3768\ : std_logic;
signal \N__3765\ : std_logic;
signal \N__3762\ : std_logic;
signal \N__3761\ : std_logic;
signal \N__3758\ : std_logic;
signal \N__3755\ : std_logic;
signal \N__3750\ : std_logic;
signal \N__3747\ : std_logic;
signal \N__3746\ : std_logic;
signal \N__3741\ : std_logic;
signal \N__3738\ : std_logic;
signal \N__3737\ : std_logic;
signal \N__3734\ : std_logic;
signal \N__3729\ : std_logic;
signal \N__3726\ : std_logic;
signal \N__3725\ : std_logic;
signal \N__3720\ : std_logic;
signal \N__3717\ : std_logic;
signal \N__3716\ : std_logic;
signal \N__3713\ : std_logic;
signal \N__3710\ : std_logic;
signal \N__3707\ : std_logic;
signal \N__3702\ : std_logic;
signal \N__3701\ : std_logic;
signal \N__3698\ : std_logic;
signal \N__3695\ : std_logic;
signal \N__3694\ : std_logic;
signal \N__3693\ : std_logic;
signal \N__3692\ : std_logic;
signal \N__3691\ : std_logic;
signal \N__3690\ : std_logic;
signal \N__3685\ : std_logic;
signal \N__3684\ : std_logic;
signal \N__3683\ : std_logic;
signal \N__3682\ : std_logic;
signal \N__3681\ : std_logic;
signal \N__3678\ : std_logic;
signal \N__3677\ : std_logic;
signal \N__3674\ : std_logic;
signal \N__3671\ : std_logic;
signal \N__3670\ : std_logic;
signal \N__3667\ : std_logic;
signal \N__3664\ : std_logic;
signal \N__3663\ : std_logic;
signal \N__3660\ : std_logic;
signal \N__3659\ : std_logic;
signal \N__3658\ : std_logic;
signal \N__3653\ : std_logic;
signal \N__3650\ : std_logic;
signal \N__3649\ : std_logic;
signal \N__3646\ : std_logic;
signal \N__3641\ : std_logic;
signal \N__3636\ : std_logic;
signal \N__3627\ : std_logic;
signal \N__3624\ : std_logic;
signal \N__3619\ : std_logic;
signal \N__3614\ : std_logic;
signal \N__3609\ : std_logic;
signal \N__3594\ : std_logic;
signal \N__3591\ : std_logic;
signal \N__3590\ : std_logic;
signal \N__3587\ : std_logic;
signal \N__3584\ : std_logic;
signal \N__3579\ : std_logic;
signal \N__3576\ : std_logic;
signal \N__3573\ : std_logic;
signal \N__3570\ : std_logic;
signal \N__3567\ : std_logic;
signal \N__3566\ : std_logic;
signal \N__3563\ : std_logic;
signal \N__3560\ : std_logic;
signal \N__3555\ : std_logic;
signal \N__3554\ : std_logic;
signal \N__3549\ : std_logic;
signal \N__3546\ : std_logic;
signal \N__3543\ : std_logic;
signal \N__3540\ : std_logic;
signal \N__3539\ : std_logic;
signal \N__3536\ : std_logic;
signal \N__3533\ : std_logic;
signal \N__3532\ : std_logic;
signal \N__3529\ : std_logic;
signal \N__3526\ : std_logic;
signal \N__3523\ : std_logic;
signal \N__3520\ : std_logic;
signal \N__3515\ : std_logic;
signal \N__3510\ : std_logic;
signal \N__3509\ : std_logic;
signal \N__3506\ : std_logic;
signal \N__3503\ : std_logic;
signal \N__3500\ : std_logic;
signal \N__3497\ : std_logic;
signal \N__3494\ : std_logic;
signal \N__3491\ : std_logic;
signal \N__3486\ : std_logic;
signal \N__3485\ : std_logic;
signal \N__3482\ : std_logic;
signal \N__3479\ : std_logic;
signal \N__3478\ : std_logic;
signal \N__3475\ : std_logic;
signal \N__3472\ : std_logic;
signal \N__3469\ : std_logic;
signal \N__3464\ : std_logic;
signal \N__3463\ : std_logic;
signal \N__3460\ : std_logic;
signal \N__3457\ : std_logic;
signal \N__3454\ : std_logic;
signal \N__3451\ : std_logic;
signal \N__3448\ : std_logic;
signal \N__3445\ : std_logic;
signal \N__3442\ : std_logic;
signal \N__3435\ : std_logic;
signal \N__3432\ : std_logic;
signal \N__3431\ : std_logic;
signal \N__3430\ : std_logic;
signal \N__3429\ : std_logic;
signal \N__3428\ : std_logic;
signal \N__3425\ : std_logic;
signal \N__3422\ : std_logic;
signal \N__3417\ : std_logic;
signal \N__3414\ : std_logic;
signal \N__3405\ : std_logic;
signal \N__3404\ : std_logic;
signal \N__3401\ : std_logic;
signal \N__3398\ : std_logic;
signal \N__3397\ : std_logic;
signal \N__3396\ : std_logic;
signal \N__3393\ : std_logic;
signal \N__3390\ : std_logic;
signal \N__3387\ : std_logic;
signal \N__3384\ : std_logic;
signal \N__3375\ : std_logic;
signal \N__3372\ : std_logic;
signal \N__3371\ : std_logic;
signal \N__3368\ : std_logic;
signal \N__3365\ : std_logic;
signal \N__3360\ : std_logic;
signal \N__3359\ : std_logic;
signal \N__3356\ : std_logic;
signal \N__3353\ : std_logic;
signal \N__3352\ : std_logic;
signal \N__3347\ : std_logic;
signal \N__3344\ : std_logic;
signal \N__3339\ : std_logic;
signal \N__3336\ : std_logic;
signal \N__3335\ : std_logic;
signal \N__3334\ : std_logic;
signal \N__3331\ : std_logic;
signal \N__3326\ : std_logic;
signal \N__3321\ : std_logic;
signal \N__3318\ : std_logic;
signal \N__3315\ : std_logic;
signal \N__3312\ : std_logic;
signal \N__3311\ : std_logic;
signal \N__3308\ : std_logic;
signal \N__3305\ : std_logic;
signal \N__3300\ : std_logic;
signal \N__3299\ : std_logic;
signal \N__3296\ : std_logic;
signal \N__3293\ : std_logic;
signal \N__3292\ : std_logic;
signal \N__3291\ : std_logic;
signal \N__3288\ : std_logic;
signal \N__3285\ : std_logic;
signal \N__3280\ : std_logic;
signal \N__3273\ : std_logic;
signal \N__3270\ : std_logic;
signal \N__3267\ : std_logic;
signal \N__3264\ : std_logic;
signal \N__3263\ : std_logic;
signal \N__3260\ : std_logic;
signal \N__3257\ : std_logic;
signal \N__3252\ : std_logic;
signal \N__3251\ : std_logic;
signal \N__3248\ : std_logic;
signal \N__3247\ : std_logic;
signal \N__3244\ : std_logic;
signal \N__3243\ : std_logic;
signal \N__3240\ : std_logic;
signal \N__3237\ : std_logic;
signal \N__3232\ : std_logic;
signal \N__3225\ : std_logic;
signal \N__3222\ : std_logic;
signal \N__3219\ : std_logic;
signal \N__3218\ : std_logic;
signal \N__3215\ : std_logic;
signal \N__3212\ : std_logic;
signal \N__3207\ : std_logic;
signal \N__3204\ : std_logic;
signal \N__3203\ : std_logic;
signal \N__3200\ : std_logic;
signal \N__3197\ : std_logic;
signal \N__3192\ : std_logic;
signal \N__3189\ : std_logic;
signal \N__3188\ : std_logic;
signal \N__3187\ : std_logic;
signal \N__3186\ : std_logic;
signal \N__3183\ : std_logic;
signal \N__3176\ : std_logic;
signal \N__3171\ : std_logic;
signal \N__3168\ : std_logic;
signal \N__3165\ : std_logic;
signal \N__3164\ : std_logic;
signal \N__3161\ : std_logic;
signal \N__3158\ : std_logic;
signal \N__3153\ : std_logic;
signal \N__3150\ : std_logic;
signal \N__3147\ : std_logic;
signal \N__3146\ : std_logic;
signal \N__3143\ : std_logic;
signal \N__3140\ : std_logic;
signal \N__3135\ : std_logic;
signal \N__3132\ : std_logic;
signal \N__3129\ : std_logic;
signal \N__3128\ : std_logic;
signal \N__3127\ : std_logic;
signal \N__3126\ : std_logic;
signal \N__3125\ : std_logic;
signal \N__3122\ : std_logic;
signal \N__3119\ : std_logic;
signal \N__3116\ : std_logic;
signal \N__3113\ : std_logic;
signal \N__3110\ : std_logic;
signal \N__3099\ : std_logic;
signal \N__3096\ : std_logic;
signal \N__3093\ : std_logic;
signal \N__3092\ : std_logic;
signal \N__3089\ : std_logic;
signal \N__3086\ : std_logic;
signal \N__3081\ : std_logic;
signal \N__3078\ : std_logic;
signal \N__3075\ : std_logic;
signal \N__3074\ : std_logic;
signal \N__3069\ : std_logic;
signal \N__3066\ : std_logic;
signal \N__3065\ : std_logic;
signal \N__3060\ : std_logic;
signal \N__3057\ : std_logic;
signal \N__3056\ : std_logic;
signal \N__3053\ : std_logic;
signal \N__3050\ : std_logic;
signal \N__3045\ : std_logic;
signal \N__3044\ : std_logic;
signal \N__3041\ : std_logic;
signal \N__3038\ : std_logic;
signal \N__3033\ : std_logic;
signal \N__3032\ : std_logic;
signal \N__3029\ : std_logic;
signal \N__3026\ : std_logic;
signal \N__3023\ : std_logic;
signal \N__3018\ : std_logic;
signal \N__3017\ : std_logic;
signal \N__3014\ : std_logic;
signal \N__3011\ : std_logic;
signal \N__3006\ : std_logic;
signal \N__3005\ : std_logic;
signal \N__3002\ : std_logic;
signal \N__2999\ : std_logic;
signal \N__2994\ : std_logic;
signal \N__2993\ : std_logic;
signal \N__2990\ : std_logic;
signal \N__2987\ : std_logic;
signal \N__2982\ : std_logic;
signal \N__2981\ : std_logic;
signal \N__2978\ : std_logic;
signal \N__2975\ : std_logic;
signal \N__2972\ : std_logic;
signal \N__2967\ : std_logic;
signal \N__2966\ : std_logic;
signal \N__2963\ : std_logic;
signal \N__2960\ : std_logic;
signal \N__2955\ : std_logic;
signal \N__2952\ : std_logic;
signal \N__2949\ : std_logic;
signal \N__2946\ : std_logic;
signal \N__2943\ : std_logic;
signal \N__2940\ : std_logic;
signal \N__2939\ : std_logic;
signal \N__2936\ : std_logic;
signal \N__2933\ : std_logic;
signal \N__2928\ : std_logic;
signal \N__2925\ : std_logic;
signal \N__2922\ : std_logic;
signal \N__2919\ : std_logic;
signal \N__2916\ : std_logic;
signal \N__2913\ : std_logic;
signal \N__2910\ : std_logic;
signal \N__2909\ : std_logic;
signal \N__2908\ : std_logic;
signal \N__2907\ : std_logic;
signal \N__2906\ : std_logic;
signal \N__2905\ : std_logic;
signal \N__2904\ : std_logic;
signal \N__2903\ : std_logic;
signal \N__2902\ : std_logic;
signal \N__2901\ : std_logic;
signal \N__2900\ : std_logic;
signal \N__2899\ : std_logic;
signal \N__2890\ : std_logic;
signal \N__2881\ : std_logic;
signal \N__2880\ : std_logic;
signal \N__2879\ : std_logic;
signal \N__2878\ : std_logic;
signal \N__2877\ : std_logic;
signal \N__2876\ : std_logic;
signal \N__2875\ : std_logic;
signal \N__2874\ : std_logic;
signal \N__2873\ : std_logic;
signal \N__2872\ : std_logic;
signal \N__2871\ : std_logic;
signal \N__2870\ : std_logic;
signal \N__2861\ : std_logic;
signal \N__2858\ : std_logic;
signal \N__2855\ : std_logic;
signal \N__2846\ : std_logic;
signal \N__2839\ : std_logic;
signal \N__2830\ : std_logic;
signal \N__2817\ : std_logic;
signal \N__2816\ : std_logic;
signal \N__2813\ : std_logic;
signal \N__2810\ : std_logic;
signal \N__2805\ : std_logic;
signal \N__2804\ : std_logic;
signal \N__2801\ : std_logic;
signal \N__2798\ : std_logic;
signal \N__2793\ : std_logic;
signal \N__2792\ : std_logic;
signal \N__2789\ : std_logic;
signal \N__2786\ : std_logic;
signal \N__2783\ : std_logic;
signal \N__2778\ : std_logic;
signal \N__2777\ : std_logic;
signal \N__2774\ : std_logic;
signal \N__2771\ : std_logic;
signal \N__2766\ : std_logic;
signal \N__2763\ : std_logic;
signal \N__2760\ : std_logic;
signal \N__2757\ : std_logic;
signal \N__2754\ : std_logic;
signal \N__2753\ : std_logic;
signal \N__2752\ : std_logic;
signal \N__2751\ : std_logic;
signal \N__2750\ : std_logic;
signal \N__2749\ : std_logic;
signal \N__2748\ : std_logic;
signal \N__2737\ : std_logic;
signal \N__2734\ : std_logic;
signal \N__2731\ : std_logic;
signal \N__2724\ : std_logic;
signal \N__2723\ : std_logic;
signal \N__2722\ : std_logic;
signal \N__2721\ : std_logic;
signal \N__2712\ : std_logic;
signal \N__2709\ : std_logic;
signal \N__2706\ : std_logic;
signal \N__2703\ : std_logic;
signal \N__2702\ : std_logic;
signal \N__2699\ : std_logic;
signal \N__2696\ : std_logic;
signal \N__2691\ : std_logic;
signal \N__2690\ : std_logic;
signal \N__2687\ : std_logic;
signal \N__2684\ : std_logic;
signal \N__2679\ : std_logic;
signal \N__2678\ : std_logic;
signal \N__2675\ : std_logic;
signal \N__2672\ : std_logic;
signal \N__2669\ : std_logic;
signal \N__2664\ : std_logic;
signal \N__2663\ : std_logic;
signal \N__2660\ : std_logic;
signal \N__2657\ : std_logic;
signal \N__2652\ : std_logic;
signal \N__2651\ : std_logic;
signal \N__2648\ : std_logic;
signal \N__2645\ : std_logic;
signal \N__2640\ : std_logic;
signal \N__2639\ : std_logic;
signal \N__2636\ : std_logic;
signal \N__2633\ : std_logic;
signal \N__2630\ : std_logic;
signal \N__2625\ : std_logic;
signal \N__2624\ : std_logic;
signal \N__2621\ : std_logic;
signal \N__2618\ : std_logic;
signal \N__2615\ : std_logic;
signal \N__2610\ : std_logic;
signal \N__2609\ : std_logic;
signal \N__2606\ : std_logic;
signal \N__2603\ : std_logic;
signal \N__2598\ : std_logic;
signal \N__2597\ : std_logic;
signal \N__2594\ : std_logic;
signal \N__2591\ : std_logic;
signal \N__2588\ : std_logic;
signal \N__2583\ : std_logic;
signal \N__2582\ : std_logic;
signal \N__2579\ : std_logic;
signal \N__2576\ : std_logic;
signal \N__2571\ : std_logic;
signal \N__2570\ : std_logic;
signal \N__2567\ : std_logic;
signal \N__2564\ : std_logic;
signal \N__2561\ : std_logic;
signal \N__2556\ : std_logic;
signal \N__2555\ : std_logic;
signal \N__2552\ : std_logic;
signal \N__2549\ : std_logic;
signal \N__2546\ : std_logic;
signal \N__2541\ : std_logic;
signal \N__2540\ : std_logic;
signal \N__2537\ : std_logic;
signal \N__2532\ : std_logic;
signal \N__2529\ : std_logic;
signal \N__2528\ : std_logic;
signal \N__2525\ : std_logic;
signal \N__2522\ : std_logic;
signal \N__2519\ : std_logic;
signal \N__2514\ : std_logic;
signal \N__2513\ : std_logic;
signal \N__2512\ : std_logic;
signal \N__2511\ : std_logic;
signal \N__2510\ : std_logic;
signal \N__2509\ : std_logic;
signal \N__2508\ : std_logic;
signal \N__2497\ : std_logic;
signal \N__2492\ : std_logic;
signal \N__2487\ : std_logic;
signal \N__2486\ : std_logic;
signal \N__2483\ : std_logic;
signal \N__2480\ : std_logic;
signal \N__2477\ : std_logic;
signal \N__2472\ : std_logic;
signal \N__2469\ : std_logic;
signal \N__2466\ : std_logic;
signal \N__2463\ : std_logic;
signal \N__2460\ : std_logic;
signal \N__2457\ : std_logic;
signal \N__2456\ : std_logic;
signal \N__2453\ : std_logic;
signal \N__2450\ : std_logic;
signal \N__2445\ : std_logic;
signal \N__2442\ : std_logic;
signal \N__2439\ : std_logic;
signal \N__2438\ : std_logic;
signal \N__2435\ : std_logic;
signal \N__2432\ : std_logic;
signal \N__2427\ : std_logic;
signal \N__2424\ : std_logic;
signal \N__2423\ : std_logic;
signal \N__2420\ : std_logic;
signal \N__2417\ : std_logic;
signal \N__2412\ : std_logic;
signal \N__2411\ : std_logic;
signal \N__2406\ : std_logic;
signal \N__2403\ : std_logic;
signal \N__2400\ : std_logic;
signal \N__2399\ : std_logic;
signal \N__2394\ : std_logic;
signal \N__2391\ : std_logic;
signal \N__2388\ : std_logic;
signal \N__2385\ : std_logic;
signal \N__2382\ : std_logic;
signal \N__2381\ : std_logic;
signal \N__2378\ : std_logic;
signal \N__2375\ : std_logic;
signal \N__2372\ : std_logic;
signal \N__2369\ : std_logic;
signal \N__2364\ : std_logic;
signal \N__2363\ : std_logic;
signal \N__2360\ : std_logic;
signal \N__2357\ : std_logic;
signal \N__2354\ : std_logic;
signal \N__2349\ : std_logic;
signal \N__2348\ : std_logic;
signal \N__2345\ : std_logic;
signal \N__2342\ : std_logic;
signal \N__2339\ : std_logic;
signal \N__2334\ : std_logic;
signal \N__2331\ : std_logic;
signal \N__2330\ : std_logic;
signal \N__2325\ : std_logic;
signal \N__2322\ : std_logic;
signal \N__2319\ : std_logic;
signal \N__2318\ : std_logic;
signal \N__2313\ : std_logic;
signal \N__2310\ : std_logic;
signal \N__2307\ : std_logic;
signal \N__2306\ : std_logic;
signal \N__2301\ : std_logic;
signal \N__2298\ : std_logic;
signal \N__2295\ : std_logic;
signal \N__2292\ : std_logic;
signal \N__2289\ : std_logic;
signal \N__2286\ : std_logic;
signal \N__2283\ : std_logic;
signal \N__2280\ : std_logic;
signal \N__2277\ : std_logic;
signal \N__2274\ : std_logic;
signal \N__2271\ : std_logic;
signal \N__2270\ : std_logic;
signal \N__2269\ : std_logic;
signal \N__2268\ : std_logic;
signal \N__2267\ : std_logic;
signal \N__2266\ : std_logic;
signal \N__2265\ : std_logic;
signal \N__2264\ : std_logic;
signal \N__2261\ : std_logic;
signal \N__2256\ : std_logic;
signal \N__2245\ : std_logic;
signal \N__2238\ : std_logic;
signal \N__2235\ : std_logic;
signal \N__2232\ : std_logic;
signal \N__2229\ : std_logic;
signal \N__2226\ : std_logic;
signal \N__2223\ : std_logic;
signal \N__2220\ : std_logic;
signal \N__2217\ : std_logic;
signal \N__2214\ : std_logic;
signal \N__2211\ : std_logic;
signal \N__2208\ : std_logic;
signal \N__2205\ : std_logic;
signal \N__2202\ : std_logic;
signal \N__2199\ : std_logic;
signal \N__2196\ : std_logic;
signal \N__2193\ : std_logic;
signal \N__2190\ : std_logic;
signal \N__2187\ : std_logic;
signal \N__2184\ : std_logic;
signal \N__2181\ : std_logic;
signal \N__2178\ : std_logic;
signal \N__2177\ : std_logic;
signal \N__2174\ : std_logic;
signal \N__2171\ : std_logic;
signal \N__2166\ : std_logic;
signal \N__2163\ : std_logic;
signal \N__2160\ : std_logic;
signal \N__2157\ : std_logic;
signal \N__2154\ : std_logic;
signal \N__2151\ : std_logic;
signal \N__2148\ : std_logic;
signal \N__2145\ : std_logic;
signal \N__2142\ : std_logic;
signal \N__2139\ : std_logic;
signal \N__2136\ : std_logic;
signal \N__2133\ : std_logic;
signal \N__2130\ : std_logic;
signal \N__2127\ : std_logic;
signal \N__2124\ : std_logic;
signal \N__2121\ : std_logic;
signal \N__2118\ : std_logic;
signal \N__2115\ : std_logic;
signal \N__2112\ : std_logic;
signal \N__2109\ : std_logic;
signal \N__2106\ : std_logic;
signal \N__2103\ : std_logic;
signal \N__2100\ : std_logic;
signal \N__2097\ : std_logic;
signal \N__2094\ : std_logic;
signal \N__2091\ : std_logic;
signal \N__2088\ : std_logic;
signal \N__2085\ : std_logic;
signal \N__2082\ : std_logic;
signal \N__2079\ : std_logic;
signal \N__2076\ : std_logic;
signal \N__2075\ : std_logic;
signal \N__2072\ : std_logic;
signal \N__2067\ : std_logic;
signal \N__2064\ : std_logic;
signal \N__2063\ : std_logic;
signal \N__2060\ : std_logic;
signal \N__2057\ : std_logic;
signal \N__2054\ : std_logic;
signal \N__2049\ : std_logic;
signal \N__2048\ : std_logic;
signal \N__2043\ : std_logic;
signal \N__2040\ : std_logic;
signal \N__2037\ : std_logic;
signal \N__2034\ : std_logic;
signal \N__2031\ : std_logic;
signal \N__2028\ : std_logic;
signal \N__2025\ : std_logic;
signal \N__2022\ : std_logic;
signal \N__2019\ : std_logic;
signal \N__2018\ : std_logic;
signal \N__2013\ : std_logic;
signal \N__2010\ : std_logic;
signal \N__2007\ : std_logic;
signal \N__2004\ : std_logic;
signal \N__2001\ : std_logic;
signal \N__1998\ : std_logic;
signal \N__1995\ : std_logic;
signal \N__1992\ : std_logic;
signal \N__1989\ : std_logic;
signal \N__1986\ : std_logic;
signal io_jtag_tck_pad_gb_input : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \n12_cascade_\ : std_logic;
signal n1307 : std_logic;
signal \n2116_cascade_\ : std_logic;
signal \n9_adj_2_cascade_\ : std_logic;
signal n8 : std_logic;
signal n12 : std_logic;
signal \n2_cascade_\ : std_logic;
signal \ctrl_idcodeArea_shifter_2\ : std_logic;
signal n1828 : std_logic;
signal \n2045_cascade_\ : std_logic;
signal \ctrl_idcodeArea_shifter_4\ : std_logic;
signal \ctrl_idcodeArea_shifter_3\ : std_logic;
signal \ctrl_idcodeArea_shifter_30\ : std_logic;
signal \n1854_cascade_\ : std_logic;
signal \n2188_cascade_\ : std_logic;
signal \n2235_cascade_\ : std_logic;
signal \n2202_cascade_\ : std_logic;
signal n2211 : std_logic;
signal n962 : std_logic;
signal n1025 : std_logic;
signal \n1025_cascade_\ : std_logic;
signal \n960_cascade_\ : std_logic;
signal n2194 : std_logic;
signal n1023 : std_logic;
signal n1027 : std_logic;
signal n965 : std_logic;
signal n5 : std_logic;
signal \n5_cascade_\ : std_logic;
signal n2201 : std_logic;
signal \bfn_1_6_0_\ : std_logic;
signal n2009 : std_logic;
signal n2010 : std_logic;
signal n2011 : std_logic;
signal n2012 : std_logic;
signal n2013 : std_logic;
signal n2014 : std_logic;
signal n2015 : std_logic;
signal n2016 : std_logic;
signal \bfn_1_7_0_\ : std_logic;
signal n2017 : std_logic;
signal n2018 : std_logic;
signal n2019 : std_logic;
signal n2020 : std_logic;
signal n2021 : std_logic;
signal n2022 : std_logic;
signal n2023 : std_logic;
signal n2024 : std_logic;
signal \bfn_1_8_0_\ : std_logic;
signal n2025 : std_logic;
signal n2026 : std_logic;
signal n2027 : std_logic;
signal n2028 : std_logic;
signal n2029 : std_logic;
signal n2030 : std_logic;
signal n2116 : std_logic;
signal \n4_cascade_\ : std_logic;
signal \ctrl_tap_tdoUnbufferd_N_223_cascade_\ : std_logic;
signal \ctrl_tap_tdoUnbufferd\ : std_logic;
signal n2146 : std_logic;
signal \n1313_cascade_\ : std_logic;
signal \ctrl_tap_tdoUnbufferd_N_224\ : std_logic;
signal \ctrl_idcodeArea_shifter_1\ : std_logic;
signal \ctrl_idcodeArea_shifter_0\ : std_logic;
signal \ctrl_idcodeArea_shifter_29\ : std_logic;
signal \ctrl_idcodeArea_shifter_28\ : std_logic;
signal \ctrl_idcodeArea_shifter_27\ : std_logic;
signal \ctrl_idcodeArea_shifter_26\ : std_logic;
signal \ctrl_idcodeArea_shifter_25\ : std_logic;
signal n6 : std_logic;
signal n1293 : std_logic;
signal \n1582_cascade_\ : std_logic;
signal n2119 : std_logic;
signal \ctrl_idcodeArea_shifter_24\ : std_logic;
signal \n2178_cascade_\ : std_logic;
signal \ctrl_idcodeArea_shifter_23\ : std_logic;
signal \ctrl_idcodeArea_shifter_5\ : std_logic;
signal \ctrl_idcodeArea_shifter_7\ : std_logic;
signal \ctrl_idcodeArea_shifter_6\ : std_logic;
signal n2045 : std_logic;
signal \ctrl_idcodeArea_shifter_8\ : std_logic;
signal n2140 : std_logic;
signal \n9_cascade_\ : std_logic;
signal n2191 : std_logic;
signal n12_adj_3 : std_logic;
signal n1769 : std_logic;
signal n1864 : std_logic;
signal \myClockArea_timeout_counter_value_3\ : std_logic;
signal \myClockArea_timeout_counter_value_1\ : std_logic;
signal \myClockArea_timeout_counter_value_5\ : std_logic;
signal \myClockArea_timeout_counter_value_0\ : std_logic;
signal \myClockArea_timeout_counter_value_9\ : std_logic;
signal \myClockArea_timeout_counter_value_18\ : std_logic;
signal \myClockArea_timeout_counter_value_12\ : std_logic;
signal \myClockArea_timeout_counter_value_14\ : std_logic;
signal \ctrl_idcodeArea_shifter_9\ : std_logic;
signal \myClockArea_timeout_counter_value_7\ : std_logic;
signal \myClockArea_timeout_counter_value_21\ : std_logic;
signal \ctrl_idcodeArea_shifter_11\ : std_logic;
signal \ctrl_idcodeArea_shifter_10\ : std_logic;
signal \myClockArea_timeout_counter_value_4\ : std_logic;
signal \myClockArea_timeout_counter_value_6\ : std_logic;
signal \myClockArea_timeout_counter_value_22\ : std_logic;
signal \myClockArea_timeout_counter_value_16\ : std_logic;
signal \myClockArea_timeout_counter_value_17\ : std_logic;
signal \myClockArea_timeout_counter_value_8\ : std_logic;
signal \myClockArea_timeout_counter_value_10\ : std_logic;
signal \myClockArea_timeout_counter_value_2\ : std_logic;
signal n2176 : std_logic;
signal \n2160_cascade_\ : std_logic;
signal n2164 : std_logic;
signal \myClockArea_timeout_counter_value_13\ : std_logic;
signal n11 : std_logic;
signal \n2182_cascade_\ : std_logic;
signal n13 : std_logic;
signal \n2113_cascade_\ : std_logic;
signal n1771 : std_logic;
signal \myClockArea_timeout_counter_value_19\ : std_logic;
signal \myClockArea_timeout_counter_value_15\ : std_logic;
signal \myClockArea_timeout_counter_value_20\ : std_logic;
signal \myClockArea_timeout_counter_value_11\ : std_logic;
signal n2162 : std_logic;
signal n2113 : std_logic;
signal global_reset_c : std_logic;
signal ctrl_tap_instruction_1 : std_logic;
signal ctrl_tap_instruction_2 : std_logic;
signal \ctrl_tap_instructionShift_2\ : std_logic;
signal ctrl_tap_instruction_4 : std_logic;
signal ctrl_tap_instruction_5 : std_logic;
signal \ctrl_tap_instructionShift_5\ : std_logic;
signal ctrl_tap_instruction_7 : std_logic;
signal \ctrl_tap_instructionShift_4\ : std_logic;
signal ctrl_tap_instruction_3 : std_logic;
signal \ctrl_tap_instructionShift_3\ : std_logic;
signal \ctrl_tap_instructionShift_7\ : std_logic;
signal ctrl_tap_instruction_6 : std_logic;
signal \ctrl_tap_instructionShift_6\ : std_logic;
signal \ctrl_tap_instructionShift_1\ : std_logic;
signal ctrl_tap_instruction_0 : std_logic;
signal \ctrl_tap_instructionShift_0\ : std_logic;
signal n15 : std_logic;
signal \ctrl_idcodeArea_shifter_18\ : std_logic;
signal \ctrl_idcodeArea_shifter_20\ : std_logic;
signal \ctrl_idcodeArea_shifter_19\ : std_logic;
signal \ctrl_idcodeArea_shifter_31\ : std_logic;
signal ctrl_tap_fsm_state_2 : std_logic;
signal n1067 : std_logic;
signal \ctrl_idcodeArea_shifter_22\ : std_logic;
signal \ctrl_idcodeArea_shifter_21\ : std_logic;
signal io_leds_c_0 : std_logic;
signal \ctrl_ledsArea_shifter_0\ : std_logic;
signal io_leds_c_1 : std_logic;
signal \ctrl_ledsArea_shifter_1\ : std_logic;
signal io_leds_c_2 : std_logic;
signal \ctrl_ledsArea_shifter_2\ : std_logic;
signal io_leds_c_3 : std_logic;
signal \ctrl_ledsArea_shifter_3\ : std_logic;
signal \ctrl_ledsArea_store_4\ : std_logic;
signal \ctrl_ledsArea_shifter_4\ : std_logic;
signal io_leds_c_5 : std_logic;
signal \ctrl_ledsArea_shifter_5\ : std_logic;
signal io_leds_c_6 : std_logic;
signal \ctrl_ledsArea_shifter_6\ : std_logic;
signal n7_adj_1 : std_logic;
signal io_leds_c_7 : std_logic;
signal n7 : std_logic;
signal \ctrl_ledsArea_shifter_7\ : std_logic;
signal n1353 : std_logic;
signal ctrl_tap_fsm_state_0 : std_logic;
signal ctrl_tap_fsm_state_3 : std_logic;
signal \ctrl_tap_fsm_stateNext_3__N_10_c_3\ : std_logic;
signal ctrl_tap_fsm_state_1 : std_logic;
signal n963 : std_logic;
signal \myClockArea_timeout_state\ : std_logic;
signal io_leds_c_4 : std_logic;
signal global_clk_c : std_logic;
signal io_jtag_tdi_c : std_logic;
signal ctrl_tap_bypass : std_logic;
signal \ctrl_idcodeArea_shifter_17\ : std_logic;
signal \ctrl_idcodeArea_shifter_14\ : std_logic;
signal \ctrl_idcodeArea_shifter_13\ : std_logic;
signal \ctrl_idcodeArea_shifter_12\ : std_logic;
signal \ctrl_idcodeArea_shifter_16\ : std_logic;
signal n2178 : std_logic;
signal n1582 : std_logic;
signal \ctrl_idcodeArea_shifter_15\ : std_logic;
signal io_jtag_tck_c : std_logic;
signal \_gnd_net_\ : std_logic;

signal global_clk_wire : std_logic;
signal io_jtag_tms_wire : std_logic;
signal global_reset_wire : std_logic;
signal io_jtag_tdi_wire : std_logic;
signal io_jtag_tdo_wire : std_logic;
signal io_leds_wire : std_logic_vector(7 downto 0);
signal io_jtag_tck_wire : std_logic;

begin
    global_clk_wire <= global_clk;
    io_jtag_tms_wire <= io_jtag_tms;
    global_reset_wire <= global_reset;
    io_jtag_tdi_wire <= io_jtag_tdi;
    io_jtag_tdo <= io_jtag_tdo_wire;
    io_leds <= io_leds_wire;
    io_jtag_tck_wire <= io_jtag_tck;

    \global_clk_pad_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__5398\,
            GLOBALBUFFEROUTPUT => global_clk_c
        );

    \global_clk_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5400\,
            DIN => \N__5399\,
            DOUT => \N__5398\,
            PACKAGEPIN => global_clk_wire
        );

    \global_clk_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__5400\,
            PADOUT => \N__5399\,
            PADIN => \N__5398\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \ctrl_tap_fsm_stateNext_3__N_10_pad_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5389\,
            DIN => \N__5388\,
            DOUT => \N__5387\,
            PACKAGEPIN => io_jtag_tms_wire
        );

    \ctrl_tap_fsm_stateNext_3__N_10_pad_3_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__5389\,
            PADOUT => \N__5388\,
            PADIN => \N__5387\,
            CLOCKENABLE => 'H',
            DIN0 => \ctrl_tap_fsm_stateNext_3__N_10_c_3\,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \global_reset_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5380\,
            DIN => \N__5379\,
            DOUT => \N__5378\,
            PACKAGEPIN => global_reset_wire
        );

    \global_reset_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__5380\,
            PADOUT => \N__5379\,
            PADIN => \N__5378\,
            CLOCKENABLE => 'H',
            DIN0 => global_reset_c,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \io_jtag_tdi_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5371\,
            DIN => \N__5370\,
            DOUT => \N__5369\,
            PACKAGEPIN => io_jtag_tdi_wire
        );

    \io_jtag_tdi_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__5371\,
            PADOUT => \N__5370\,
            PADIN => \N__5369\,
            CLOCKENABLE => 'H',
            DIN0 => io_jtag_tdi_c,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \io_jtag_tdo_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5362\,
            DIN => \N__5361\,
            DOUT => \N__5360\,
            PACKAGEPIN => io_jtag_tdo_wire
        );

    \io_jtag_tdo_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "010101",
            NEG_TRIGGER => '1'
        )
    port map (
            PADOEN => \N__5362\,
            PADOUT => \N__5361\,
            PADIN => \N__5360\,
            CLOCKENABLE => \VCCG0\,
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__2283\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => \N__4716\,
            OUTPUTENABLE => '0'
        );

    \io_leds_pad_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5353\,
            DIN => \N__5352\,
            DOUT => \N__5351\,
            PACKAGEPIN => io_leds_wire(0)
        );

    \io_leds_pad_0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__5353\,
            PADOUT => \N__5352\,
            PADIN => \N__5351\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__3546\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \io_leds_pad_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5344\,
            DIN => \N__5343\,
            DOUT => \N__5342\,
            PACKAGEPIN => io_leds_wire(1)
        );

    \io_leds_pad_1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__5344\,
            PADOUT => \N__5343\,
            PADIN => \N__5342\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__4659\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \io_leds_pad_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5335\,
            DIN => \N__5334\,
            DOUT => \N__5333\,
            PACKAGEPIN => io_leds_wire(2)
        );

    \io_leds_pad_2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__5335\,
            PADOUT => \N__5334\,
            PADIN => \N__5333\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__4605\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \io_leds_pad_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5326\,
            DIN => \N__5325\,
            DOUT => \N__5324\,
            PACKAGEPIN => io_leds_wire(3)
        );

    \io_leds_pad_3_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__5326\,
            PADOUT => \N__5325\,
            PADIN => \N__5324\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__4557\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \io_leds_pad_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5317\,
            DIN => \N__5316\,
            DOUT => \N__5315\,
            PACKAGEPIN => io_leds_wire(4)
        );

    \io_leds_pad_4_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__5317\,
            PADOUT => \N__5316\,
            PADIN => \N__5315\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__5238\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \io_leds_pad_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5308\,
            DIN => \N__5307\,
            DOUT => \N__5306\,
            PACKAGEPIN => io_leds_wire(5)
        );

    \io_leds_pad_5_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__5308\,
            PADOUT => \N__5307\,
            PADIN => \N__5306\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__4464\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \io_leds_pad_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5299\,
            DIN => \N__5298\,
            DOUT => \N__5297\,
            PACKAGEPIN => io_leds_wire(6)
        );

    \io_leds_pad_6_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__5299\,
            PADOUT => \N__5298\,
            PADIN => \N__5297\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__4412\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \io_leds_pad_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5290\,
            DIN => \N__5289\,
            DOUT => \N__5288\,
            PACKAGEPIN => io_leds_wire(7)
        );

    \io_leds_pad_7_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__5290\,
            PADOUT => \N__5289\,
            PADIN => \N__5288\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__4320\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \io_jtag_tck_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5281\,
            DIN => \N__5280\,
            DOUT => \N__5279\,
            PACKAGEPIN => io_jtag_tck_wire
        );

    \io_jtag_tck_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__5281\,
            PADOUT => \N__5280\,
            PADIN => \N__5279\,
            CLOCKENABLE => 'H',
            DIN0 => io_jtag_tck_pad_gb_input,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \I__1261\ : InMux
    port map (
            O => \N__5262\,
            I => \N__5258\
        );

    \I__1260\ : InMux
    port map (
            O => \N__5261\,
            I => \N__5254\
        );

    \I__1259\ : LocalMux
    port map (
            O => \N__5258\,
            I => \N__5251\
        );

    \I__1258\ : InMux
    port map (
            O => \N__5257\,
            I => \N__5248\
        );

    \I__1257\ : LocalMux
    port map (
            O => \N__5254\,
            I => \N__5245\
        );

    \I__1256\ : Odrv4
    port map (
            O => \N__5251\,
            I => \myClockArea_timeout_state\
        );

    \I__1255\ : LocalMux
    port map (
            O => \N__5248\,
            I => \myClockArea_timeout_state\
        );

    \I__1254\ : Odrv4
    port map (
            O => \N__5245\,
            I => \myClockArea_timeout_state\
        );

    \I__1253\ : IoInMux
    port map (
            O => \N__5238\,
            I => \N__5235\
        );

    \I__1252\ : LocalMux
    port map (
            O => \N__5235\,
            I => \N__5232\
        );

    \I__1251\ : IoSpan4Mux
    port map (
            O => \N__5232\,
            I => \N__5229\
        );

    \I__1250\ : Sp12to4
    port map (
            O => \N__5229\,
            I => \N__5225\
        );

    \I__1249\ : InMux
    port map (
            O => \N__5228\,
            I => \N__5222\
        );

    \I__1248\ : Odrv12
    port map (
            O => \N__5225\,
            I => io_leds_c_4
        );

    \I__1247\ : LocalMux
    port map (
            O => \N__5222\,
            I => io_leds_c_4
        );

    \I__1246\ : ClkMux
    port map (
            O => \N__5217\,
            I => \N__5202\
        );

    \I__1245\ : ClkMux
    port map (
            O => \N__5216\,
            I => \N__5202\
        );

    \I__1244\ : ClkMux
    port map (
            O => \N__5215\,
            I => \N__5202\
        );

    \I__1243\ : ClkMux
    port map (
            O => \N__5214\,
            I => \N__5202\
        );

    \I__1242\ : ClkMux
    port map (
            O => \N__5213\,
            I => \N__5202\
        );

    \I__1241\ : GlobalMux
    port map (
            O => \N__5202\,
            I => \N__5199\
        );

    \I__1240\ : gio2CtrlBuf
    port map (
            O => \N__5199\,
            I => global_clk_c
        );

    \I__1239\ : CascadeMux
    port map (
            O => \N__5196\,
            I => \N__5192\
        );

    \I__1238\ : CascadeMux
    port map (
            O => \N__5195\,
            I => \N__5189\
        );

    \I__1237\ : InMux
    port map (
            O => \N__5192\,
            I => \N__5186\
        );

    \I__1236\ : InMux
    port map (
            O => \N__5189\,
            I => \N__5182\
        );

    \I__1235\ : LocalMux
    port map (
            O => \N__5186\,
            I => \N__5178\
        );

    \I__1234\ : InMux
    port map (
            O => \N__5185\,
            I => \N__5175\
        );

    \I__1233\ : LocalMux
    port map (
            O => \N__5182\,
            I => \N__5172\
        );

    \I__1232\ : InMux
    port map (
            O => \N__5181\,
            I => \N__5169\
        );

    \I__1231\ : Span4Mux_v
    port map (
            O => \N__5178\,
            I => \N__5164\
        );

    \I__1230\ : LocalMux
    port map (
            O => \N__5175\,
            I => \N__5164\
        );

    \I__1229\ : Odrv4
    port map (
            O => \N__5172\,
            I => io_jtag_tdi_c
        );

    \I__1228\ : LocalMux
    port map (
            O => \N__5169\,
            I => io_jtag_tdi_c
        );

    \I__1227\ : Odrv4
    port map (
            O => \N__5164\,
            I => io_jtag_tdi_c
        );

    \I__1226\ : InMux
    port map (
            O => \N__5157\,
            I => \N__5154\
        );

    \I__1225\ : LocalMux
    port map (
            O => \N__5154\,
            I => \N__5151\
        );

    \I__1224\ : Odrv4
    port map (
            O => \N__5151\,
            I => ctrl_tap_bypass
        );

    \I__1223\ : CascadeMux
    port map (
            O => \N__5148\,
            I => \N__5145\
        );

    \I__1222\ : InMux
    port map (
            O => \N__5145\,
            I => \N__5141\
        );

    \I__1221\ : InMux
    port map (
            O => \N__5144\,
            I => \N__5138\
        );

    \I__1220\ : LocalMux
    port map (
            O => \N__5141\,
            I => \ctrl_idcodeArea_shifter_17\
        );

    \I__1219\ : LocalMux
    port map (
            O => \N__5138\,
            I => \ctrl_idcodeArea_shifter_17\
        );

    \I__1218\ : InMux
    port map (
            O => \N__5133\,
            I => \N__5127\
        );

    \I__1217\ : InMux
    port map (
            O => \N__5132\,
            I => \N__5127\
        );

    \I__1216\ : LocalMux
    port map (
            O => \N__5127\,
            I => \ctrl_idcodeArea_shifter_14\
        );

    \I__1215\ : CascadeMux
    port map (
            O => \N__5124\,
            I => \N__5121\
        );

    \I__1214\ : InMux
    port map (
            O => \N__5121\,
            I => \N__5115\
        );

    \I__1213\ : InMux
    port map (
            O => \N__5120\,
            I => \N__5115\
        );

    \I__1212\ : LocalMux
    port map (
            O => \N__5115\,
            I => \ctrl_idcodeArea_shifter_13\
        );

    \I__1211\ : CascadeMux
    port map (
            O => \N__5112\,
            I => \N__5109\
        );

    \I__1210\ : InMux
    port map (
            O => \N__5109\,
            I => \N__5106\
        );

    \I__1209\ : LocalMux
    port map (
            O => \N__5106\,
            I => \N__5103\
        );

    \I__1208\ : Span4Mux_h
    port map (
            O => \N__5103\,
            I => \N__5099\
        );

    \I__1207\ : InMux
    port map (
            O => \N__5102\,
            I => \N__5096\
        );

    \I__1206\ : Odrv4
    port map (
            O => \N__5099\,
            I => \ctrl_idcodeArea_shifter_12\
        );

    \I__1205\ : LocalMux
    port map (
            O => \N__5096\,
            I => \ctrl_idcodeArea_shifter_12\
        );

    \I__1204\ : InMux
    port map (
            O => \N__5091\,
            I => \N__5085\
        );

    \I__1203\ : InMux
    port map (
            O => \N__5090\,
            I => \N__5085\
        );

    \I__1202\ : LocalMux
    port map (
            O => \N__5085\,
            I => \ctrl_idcodeArea_shifter_16\
        );

    \I__1201\ : CascadeMux
    port map (
            O => \N__5082\,
            I => \N__5079\
        );

    \I__1200\ : InMux
    port map (
            O => \N__5079\,
            I => \N__5071\
        );

    \I__1199\ : InMux
    port map (
            O => \N__5078\,
            I => \N__5068\
        );

    \I__1198\ : CascadeMux
    port map (
            O => \N__5077\,
            I => \N__5065\
        );

    \I__1197\ : CascadeMux
    port map (
            O => \N__5076\,
            I => \N__5058\
        );

    \I__1196\ : InMux
    port map (
            O => \N__5075\,
            I => \N__5032\
        );

    \I__1195\ : InMux
    port map (
            O => \N__5074\,
            I => \N__5032\
        );

    \I__1194\ : LocalMux
    port map (
            O => \N__5071\,
            I => \N__5027\
        );

    \I__1193\ : LocalMux
    port map (
            O => \N__5068\,
            I => \N__5027\
        );

    \I__1192\ : InMux
    port map (
            O => \N__5065\,
            I => \N__5024\
        );

    \I__1191\ : InMux
    port map (
            O => \N__5064\,
            I => \N__5021\
        );

    \I__1190\ : InMux
    port map (
            O => \N__5063\,
            I => \N__5014\
        );

    \I__1189\ : InMux
    port map (
            O => \N__5062\,
            I => \N__5014\
        );

    \I__1188\ : InMux
    port map (
            O => \N__5061\,
            I => \N__5014\
        );

    \I__1187\ : InMux
    port map (
            O => \N__5058\,
            I => \N__5011\
        );

    \I__1186\ : InMux
    port map (
            O => \N__5057\,
            I => \N__5002\
        );

    \I__1185\ : InMux
    port map (
            O => \N__5056\,
            I => \N__5002\
        );

    \I__1184\ : InMux
    port map (
            O => \N__5055\,
            I => \N__5002\
        );

    \I__1183\ : InMux
    port map (
            O => \N__5054\,
            I => \N__5002\
        );

    \I__1182\ : InMux
    port map (
            O => \N__5053\,
            I => \N__4991\
        );

    \I__1181\ : InMux
    port map (
            O => \N__5052\,
            I => \N__4991\
        );

    \I__1180\ : InMux
    port map (
            O => \N__5051\,
            I => \N__4991\
        );

    \I__1179\ : InMux
    port map (
            O => \N__5050\,
            I => \N__4991\
        );

    \I__1178\ : InMux
    port map (
            O => \N__5049\,
            I => \N__4991\
        );

    \I__1177\ : InMux
    port map (
            O => \N__5048\,
            I => \N__4986\
        );

    \I__1176\ : InMux
    port map (
            O => \N__5047\,
            I => \N__4986\
        );

    \I__1175\ : InMux
    port map (
            O => \N__5046\,
            I => \N__4979\
        );

    \I__1174\ : InMux
    port map (
            O => \N__5045\,
            I => \N__4979\
        );

    \I__1173\ : InMux
    port map (
            O => \N__5044\,
            I => \N__4979\
        );

    \I__1172\ : InMux
    port map (
            O => \N__5043\,
            I => \N__4968\
        );

    \I__1171\ : InMux
    port map (
            O => \N__5042\,
            I => \N__4968\
        );

    \I__1170\ : InMux
    port map (
            O => \N__5041\,
            I => \N__4968\
        );

    \I__1169\ : InMux
    port map (
            O => \N__5040\,
            I => \N__4968\
        );

    \I__1168\ : InMux
    port map (
            O => \N__5039\,
            I => \N__4968\
        );

    \I__1167\ : InMux
    port map (
            O => \N__5038\,
            I => \N__4963\
        );

    \I__1166\ : InMux
    port map (
            O => \N__5037\,
            I => \N__4963\
        );

    \I__1165\ : LocalMux
    port map (
            O => \N__5032\,
            I => \N__4956\
        );

    \I__1164\ : Span12Mux_s2_v
    port map (
            O => \N__5027\,
            I => \N__4956\
        );

    \I__1163\ : LocalMux
    port map (
            O => \N__5024\,
            I => \N__4956\
        );

    \I__1162\ : LocalMux
    port map (
            O => \N__5021\,
            I => \N__4951\
        );

    \I__1161\ : LocalMux
    port map (
            O => \N__5014\,
            I => \N__4951\
        );

    \I__1160\ : LocalMux
    port map (
            O => \N__5011\,
            I => \N__4944\
        );

    \I__1159\ : LocalMux
    port map (
            O => \N__5002\,
            I => \N__4944\
        );

    \I__1158\ : LocalMux
    port map (
            O => \N__4991\,
            I => \N__4944\
        );

    \I__1157\ : LocalMux
    port map (
            O => \N__4986\,
            I => n2178
        );

    \I__1156\ : LocalMux
    port map (
            O => \N__4979\,
            I => n2178
        );

    \I__1155\ : LocalMux
    port map (
            O => \N__4968\,
            I => n2178
        );

    \I__1154\ : LocalMux
    port map (
            O => \N__4963\,
            I => n2178
        );

    \I__1153\ : Odrv12
    port map (
            O => \N__4956\,
            I => n2178
        );

    \I__1152\ : Odrv4
    port map (
            O => \N__4951\,
            I => n2178
        );

    \I__1151\ : Odrv4
    port map (
            O => \N__4944\,
            I => n2178
        );

    \I__1150\ : CascadeMux
    port map (
            O => \N__4929\,
            I => \N__4907\
        );

    \I__1149\ : CascadeMux
    port map (
            O => \N__4928\,
            I => \N__4901\
        );

    \I__1148\ : InMux
    port map (
            O => \N__4927\,
            I => \N__4885\
        );

    \I__1147\ : InMux
    port map (
            O => \N__4926\,
            I => \N__4885\
        );

    \I__1146\ : InMux
    port map (
            O => \N__4925\,
            I => \N__4885\
        );

    \I__1145\ : InMux
    port map (
            O => \N__4924\,
            I => \N__4885\
        );

    \I__1144\ : InMux
    port map (
            O => \N__4923\,
            I => \N__4885\
        );

    \I__1143\ : InMux
    port map (
            O => \N__4922\,
            I => \N__4878\
        );

    \I__1142\ : InMux
    port map (
            O => \N__4921\,
            I => \N__4878\
        );

    \I__1141\ : InMux
    port map (
            O => \N__4920\,
            I => \N__4878\
        );

    \I__1140\ : CascadeMux
    port map (
            O => \N__4919\,
            I => \N__4874\
        );

    \I__1139\ : CascadeMux
    port map (
            O => \N__4918\,
            I => \N__4871\
        );

    \I__1138\ : CascadeMux
    port map (
            O => \N__4917\,
            I => \N__4867\
        );

    \I__1137\ : CascadeMux
    port map (
            O => \N__4916\,
            I => \N__4860\
        );

    \I__1136\ : InMux
    port map (
            O => \N__4915\,
            I => \N__4851\
        );

    \I__1135\ : InMux
    port map (
            O => \N__4914\,
            I => \N__4848\
        );

    \I__1134\ : InMux
    port map (
            O => \N__4913\,
            I => \N__4841\
        );

    \I__1133\ : InMux
    port map (
            O => \N__4912\,
            I => \N__4841\
        );

    \I__1132\ : InMux
    port map (
            O => \N__4911\,
            I => \N__4841\
        );

    \I__1131\ : InMux
    port map (
            O => \N__4910\,
            I => \N__4832\
        );

    \I__1130\ : InMux
    port map (
            O => \N__4907\,
            I => \N__4832\
        );

    \I__1129\ : InMux
    port map (
            O => \N__4906\,
            I => \N__4832\
        );

    \I__1128\ : InMux
    port map (
            O => \N__4905\,
            I => \N__4832\
        );

    \I__1127\ : InMux
    port map (
            O => \N__4904\,
            I => \N__4825\
        );

    \I__1126\ : InMux
    port map (
            O => \N__4901\,
            I => \N__4825\
        );

    \I__1125\ : InMux
    port map (
            O => \N__4900\,
            I => \N__4825\
        );

    \I__1124\ : InMux
    port map (
            O => \N__4899\,
            I => \N__4822\
        );

    \I__1123\ : InMux
    port map (
            O => \N__4898\,
            I => \N__4815\
        );

    \I__1122\ : InMux
    port map (
            O => \N__4897\,
            I => \N__4815\
        );

    \I__1121\ : InMux
    port map (
            O => \N__4896\,
            I => \N__4815\
        );

    \I__1120\ : LocalMux
    port map (
            O => \N__4885\,
            I => \N__4810\
        );

    \I__1119\ : LocalMux
    port map (
            O => \N__4878\,
            I => \N__4810\
        );

    \I__1118\ : InMux
    port map (
            O => \N__4877\,
            I => \N__4807\
        );

    \I__1117\ : InMux
    port map (
            O => \N__4874\,
            I => \N__4804\
        );

    \I__1116\ : InMux
    port map (
            O => \N__4871\,
            I => \N__4801\
        );

    \I__1115\ : InMux
    port map (
            O => \N__4870\,
            I => \N__4796\
        );

    \I__1114\ : InMux
    port map (
            O => \N__4867\,
            I => \N__4796\
        );

    \I__1113\ : InMux
    port map (
            O => \N__4866\,
            I => \N__4791\
        );

    \I__1112\ : InMux
    port map (
            O => \N__4865\,
            I => \N__4791\
        );

    \I__1111\ : InMux
    port map (
            O => \N__4864\,
            I => \N__4786\
        );

    \I__1110\ : InMux
    port map (
            O => \N__4863\,
            I => \N__4786\
        );

    \I__1109\ : InMux
    port map (
            O => \N__4860\,
            I => \N__4779\
        );

    \I__1108\ : InMux
    port map (
            O => \N__4859\,
            I => \N__4779\
        );

    \I__1107\ : InMux
    port map (
            O => \N__4858\,
            I => \N__4779\
        );

    \I__1106\ : InMux
    port map (
            O => \N__4857\,
            I => \N__4770\
        );

    \I__1105\ : InMux
    port map (
            O => \N__4856\,
            I => \N__4770\
        );

    \I__1104\ : InMux
    port map (
            O => \N__4855\,
            I => \N__4770\
        );

    \I__1103\ : InMux
    port map (
            O => \N__4854\,
            I => \N__4770\
        );

    \I__1102\ : LocalMux
    port map (
            O => \N__4851\,
            I => \N__4767\
        );

    \I__1101\ : LocalMux
    port map (
            O => \N__4848\,
            I => \N__4758\
        );

    \I__1100\ : LocalMux
    port map (
            O => \N__4841\,
            I => \N__4758\
        );

    \I__1099\ : LocalMux
    port map (
            O => \N__4832\,
            I => \N__4758\
        );

    \I__1098\ : LocalMux
    port map (
            O => \N__4825\,
            I => \N__4758\
        );

    \I__1097\ : LocalMux
    port map (
            O => \N__4822\,
            I => \N__4751\
        );

    \I__1096\ : LocalMux
    port map (
            O => \N__4815\,
            I => \N__4751\
        );

    \I__1095\ : Span4Mux_s1_v
    port map (
            O => \N__4810\,
            I => \N__4751\
        );

    \I__1094\ : LocalMux
    port map (
            O => \N__4807\,
            I => n1582
        );

    \I__1093\ : LocalMux
    port map (
            O => \N__4804\,
            I => n1582
        );

    \I__1092\ : LocalMux
    port map (
            O => \N__4801\,
            I => n1582
        );

    \I__1091\ : LocalMux
    port map (
            O => \N__4796\,
            I => n1582
        );

    \I__1090\ : LocalMux
    port map (
            O => \N__4791\,
            I => n1582
        );

    \I__1089\ : LocalMux
    port map (
            O => \N__4786\,
            I => n1582
        );

    \I__1088\ : LocalMux
    port map (
            O => \N__4779\,
            I => n1582
        );

    \I__1087\ : LocalMux
    port map (
            O => \N__4770\,
            I => n1582
        );

    \I__1086\ : Odrv4
    port map (
            O => \N__4767\,
            I => n1582
        );

    \I__1085\ : Odrv4
    port map (
            O => \N__4758\,
            I => n1582
        );

    \I__1084\ : Odrv4
    port map (
            O => \N__4751\,
            I => n1582
        );

    \I__1083\ : CascadeMux
    port map (
            O => \N__4728\,
            I => \N__4724\
        );

    \I__1082\ : InMux
    port map (
            O => \N__4727\,
            I => \N__4719\
        );

    \I__1081\ : InMux
    port map (
            O => \N__4724\,
            I => \N__4719\
        );

    \I__1080\ : LocalMux
    port map (
            O => \N__4719\,
            I => \ctrl_idcodeArea_shifter_15\
        );

    \I__1079\ : ClkMux
    port map (
            O => \N__4716\,
            I => \N__4665\
        );

    \I__1078\ : ClkMux
    port map (
            O => \N__4715\,
            I => \N__4665\
        );

    \I__1077\ : ClkMux
    port map (
            O => \N__4714\,
            I => \N__4665\
        );

    \I__1076\ : ClkMux
    port map (
            O => \N__4713\,
            I => \N__4665\
        );

    \I__1075\ : ClkMux
    port map (
            O => \N__4712\,
            I => \N__4665\
        );

    \I__1074\ : ClkMux
    port map (
            O => \N__4711\,
            I => \N__4665\
        );

    \I__1073\ : ClkMux
    port map (
            O => \N__4710\,
            I => \N__4665\
        );

    \I__1072\ : ClkMux
    port map (
            O => \N__4709\,
            I => \N__4665\
        );

    \I__1071\ : ClkMux
    port map (
            O => \N__4708\,
            I => \N__4665\
        );

    \I__1070\ : ClkMux
    port map (
            O => \N__4707\,
            I => \N__4665\
        );

    \I__1069\ : ClkMux
    port map (
            O => \N__4706\,
            I => \N__4665\
        );

    \I__1068\ : ClkMux
    port map (
            O => \N__4705\,
            I => \N__4665\
        );

    \I__1067\ : ClkMux
    port map (
            O => \N__4704\,
            I => \N__4665\
        );

    \I__1066\ : ClkMux
    port map (
            O => \N__4703\,
            I => \N__4665\
        );

    \I__1065\ : ClkMux
    port map (
            O => \N__4702\,
            I => \N__4665\
        );

    \I__1064\ : ClkMux
    port map (
            O => \N__4701\,
            I => \N__4665\
        );

    \I__1063\ : ClkMux
    port map (
            O => \N__4700\,
            I => \N__4665\
        );

    \I__1062\ : GlobalMux
    port map (
            O => \N__4665\,
            I => \N__4662\
        );

    \I__1061\ : gio2CtrlBuf
    port map (
            O => \N__4662\,
            I => io_jtag_tck_c
        );

    \I__1060\ : IoInMux
    port map (
            O => \N__4659\,
            I => \N__4656\
        );

    \I__1059\ : LocalMux
    port map (
            O => \N__4656\,
            I => \N__4653\
        );

    \I__1058\ : Span4Mux_s2_h
    port map (
            O => \N__4653\,
            I => \N__4650\
        );

    \I__1057\ : Span4Mux_h
    port map (
            O => \N__4650\,
            I => \N__4646\
        );

    \I__1056\ : CascadeMux
    port map (
            O => \N__4649\,
            I => \N__4643\
        );

    \I__1055\ : Span4Mux_v
    port map (
            O => \N__4646\,
            I => \N__4640\
        );

    \I__1054\ : InMux
    port map (
            O => \N__4643\,
            I => \N__4637\
        );

    \I__1053\ : Span4Mux_v
    port map (
            O => \N__4640\,
            I => \N__4631\
        );

    \I__1052\ : LocalMux
    port map (
            O => \N__4637\,
            I => \N__4631\
        );

    \I__1051\ : InMux
    port map (
            O => \N__4636\,
            I => \N__4628\
        );

    \I__1050\ : Odrv4
    port map (
            O => \N__4631\,
            I => io_leds_c_1
        );

    \I__1049\ : LocalMux
    port map (
            O => \N__4628\,
            I => io_leds_c_1
        );

    \I__1048\ : InMux
    port map (
            O => \N__4623\,
            I => \N__4619\
        );

    \I__1047\ : CascadeMux
    port map (
            O => \N__4622\,
            I => \N__4616\
        );

    \I__1046\ : LocalMux
    port map (
            O => \N__4619\,
            I => \N__4613\
        );

    \I__1045\ : InMux
    port map (
            O => \N__4616\,
            I => \N__4610\
        );

    \I__1044\ : Odrv4
    port map (
            O => \N__4613\,
            I => \ctrl_ledsArea_shifter_1\
        );

    \I__1043\ : LocalMux
    port map (
            O => \N__4610\,
            I => \ctrl_ledsArea_shifter_1\
        );

    \I__1042\ : IoInMux
    port map (
            O => \N__4605\,
            I => \N__4602\
        );

    \I__1041\ : LocalMux
    port map (
            O => \N__4602\,
            I => \N__4599\
        );

    \I__1040\ : Span4Mux_s3_h
    port map (
            O => \N__4599\,
            I => \N__4596\
        );

    \I__1039\ : Sp12to4
    port map (
            O => \N__4596\,
            I => \N__4592\
        );

    \I__1038\ : InMux
    port map (
            O => \N__4595\,
            I => \N__4589\
        );

    \I__1037\ : Span12Mux_v
    port map (
            O => \N__4592\,
            I => \N__4583\
        );

    \I__1036\ : LocalMux
    port map (
            O => \N__4589\,
            I => \N__4583\
        );

    \I__1035\ : InMux
    port map (
            O => \N__4588\,
            I => \N__4580\
        );

    \I__1034\ : Odrv12
    port map (
            O => \N__4583\,
            I => io_leds_c_2
        );

    \I__1033\ : LocalMux
    port map (
            O => \N__4580\,
            I => io_leds_c_2
        );

    \I__1032\ : InMux
    port map (
            O => \N__4575\,
            I => \N__4572\
        );

    \I__1031\ : LocalMux
    port map (
            O => \N__4572\,
            I => \N__4568\
        );

    \I__1030\ : InMux
    port map (
            O => \N__4571\,
            I => \N__4565\
        );

    \I__1029\ : Span4Mux_s2_h
    port map (
            O => \N__4568\,
            I => \N__4560\
        );

    \I__1028\ : LocalMux
    port map (
            O => \N__4565\,
            I => \N__4560\
        );

    \I__1027\ : Odrv4
    port map (
            O => \N__4560\,
            I => \ctrl_ledsArea_shifter_2\
        );

    \I__1026\ : IoInMux
    port map (
            O => \N__4557\,
            I => \N__4554\
        );

    \I__1025\ : LocalMux
    port map (
            O => \N__4554\,
            I => \N__4551\
        );

    \I__1024\ : IoSpan4Mux
    port map (
            O => \N__4551\,
            I => \N__4548\
        );

    \I__1023\ : Span4Mux_s3_h
    port map (
            O => \N__4548\,
            I => \N__4545\
        );

    \I__1022\ : Span4Mux_h
    port map (
            O => \N__4545\,
            I => \N__4541\
        );

    \I__1021\ : InMux
    port map (
            O => \N__4544\,
            I => \N__4538\
        );

    \I__1020\ : Span4Mux_v
    port map (
            O => \N__4541\,
            I => \N__4532\
        );

    \I__1019\ : LocalMux
    port map (
            O => \N__4538\,
            I => \N__4532\
        );

    \I__1018\ : InMux
    port map (
            O => \N__4537\,
            I => \N__4529\
        );

    \I__1017\ : Odrv4
    port map (
            O => \N__4532\,
            I => io_leds_c_3
        );

    \I__1016\ : LocalMux
    port map (
            O => \N__4529\,
            I => io_leds_c_3
        );

    \I__1015\ : CascadeMux
    port map (
            O => \N__4524\,
            I => \N__4521\
        );

    \I__1014\ : InMux
    port map (
            O => \N__4521\,
            I => \N__4517\
        );

    \I__1013\ : CascadeMux
    port map (
            O => \N__4520\,
            I => \N__4514\
        );

    \I__1012\ : LocalMux
    port map (
            O => \N__4517\,
            I => \N__4511\
        );

    \I__1011\ : InMux
    port map (
            O => \N__4514\,
            I => \N__4508\
        );

    \I__1010\ : Odrv4
    port map (
            O => \N__4511\,
            I => \ctrl_ledsArea_shifter_3\
        );

    \I__1009\ : LocalMux
    port map (
            O => \N__4508\,
            I => \ctrl_ledsArea_shifter_3\
        );

    \I__1008\ : InMux
    port map (
            O => \N__4503\,
            I => \N__4500\
        );

    \I__1007\ : LocalMux
    port map (
            O => \N__4500\,
            I => \N__4497\
        );

    \I__1006\ : Span4Mux_h
    port map (
            O => \N__4497\,
            I => \N__4493\
        );

    \I__1005\ : InMux
    port map (
            O => \N__4496\,
            I => \N__4490\
        );

    \I__1004\ : Odrv4
    port map (
            O => \N__4493\,
            I => \ctrl_ledsArea_store_4\
        );

    \I__1003\ : LocalMux
    port map (
            O => \N__4490\,
            I => \ctrl_ledsArea_store_4\
        );

    \I__1002\ : InMux
    port map (
            O => \N__4485\,
            I => \N__4482\
        );

    \I__1001\ : LocalMux
    port map (
            O => \N__4482\,
            I => \N__4478\
        );

    \I__1000\ : CascadeMux
    port map (
            O => \N__4481\,
            I => \N__4475\
        );

    \I__999\ : Span4Mux_s3_h
    port map (
            O => \N__4478\,
            I => \N__4472\
        );

    \I__998\ : InMux
    port map (
            O => \N__4475\,
            I => \N__4469\
        );

    \I__997\ : Odrv4
    port map (
            O => \N__4472\,
            I => \ctrl_ledsArea_shifter_4\
        );

    \I__996\ : LocalMux
    port map (
            O => \N__4469\,
            I => \ctrl_ledsArea_shifter_4\
        );

    \I__995\ : IoInMux
    port map (
            O => \N__4464\,
            I => \N__4461\
        );

    \I__994\ : LocalMux
    port map (
            O => \N__4461\,
            I => \N__4458\
        );

    \I__993\ : Span4Mux_s1_h
    port map (
            O => \N__4458\,
            I => \N__4454\
        );

    \I__992\ : InMux
    port map (
            O => \N__4457\,
            I => \N__4451\
        );

    \I__991\ : Span4Mux_v
    port map (
            O => \N__4454\,
            I => \N__4447\
        );

    \I__990\ : LocalMux
    port map (
            O => \N__4451\,
            I => \N__4444\
        );

    \I__989\ : InMux
    port map (
            O => \N__4450\,
            I => \N__4441\
        );

    \I__988\ : Odrv4
    port map (
            O => \N__4447\,
            I => io_leds_c_5
        );

    \I__987\ : Odrv12
    port map (
            O => \N__4444\,
            I => io_leds_c_5
        );

    \I__986\ : LocalMux
    port map (
            O => \N__4441\,
            I => io_leds_c_5
        );

    \I__985\ : CascadeMux
    port map (
            O => \N__4434\,
            I => \N__4431\
        );

    \I__984\ : InMux
    port map (
            O => \N__4431\,
            I => \N__4428\
        );

    \I__983\ : LocalMux
    port map (
            O => \N__4428\,
            I => \N__4424\
        );

    \I__982\ : InMux
    port map (
            O => \N__4427\,
            I => \N__4421\
        );

    \I__981\ : Odrv4
    port map (
            O => \N__4424\,
            I => \ctrl_ledsArea_shifter_5\
        );

    \I__980\ : LocalMux
    port map (
            O => \N__4421\,
            I => \ctrl_ledsArea_shifter_5\
        );

    \I__979\ : InMux
    port map (
            O => \N__4416\,
            I => \N__4413\
        );

    \I__978\ : LocalMux
    port map (
            O => \N__4413\,
            I => \N__4409\
        );

    \I__977\ : IoInMux
    port map (
            O => \N__4412\,
            I => \N__4405\
        );

    \I__976\ : Span4Mux_h
    port map (
            O => \N__4409\,
            I => \N__4402\
        );

    \I__975\ : InMux
    port map (
            O => \N__4408\,
            I => \N__4399\
        );

    \I__974\ : LocalMux
    port map (
            O => \N__4405\,
            I => io_leds_c_6
        );

    \I__973\ : Odrv4
    port map (
            O => \N__4402\,
            I => io_leds_c_6
        );

    \I__972\ : LocalMux
    port map (
            O => \N__4399\,
            I => io_leds_c_6
        );

    \I__971\ : InMux
    port map (
            O => \N__4392\,
            I => \N__4389\
        );

    \I__970\ : LocalMux
    port map (
            O => \N__4389\,
            I => \N__4385\
        );

    \I__969\ : CascadeMux
    port map (
            O => \N__4388\,
            I => \N__4382\
        );

    \I__968\ : Span4Mux_s3_h
    port map (
            O => \N__4385\,
            I => \N__4379\
        );

    \I__967\ : InMux
    port map (
            O => \N__4382\,
            I => \N__4376\
        );

    \I__966\ : Odrv4
    port map (
            O => \N__4379\,
            I => \ctrl_ledsArea_shifter_6\
        );

    \I__965\ : LocalMux
    port map (
            O => \N__4376\,
            I => \ctrl_ledsArea_shifter_6\
        );

    \I__964\ : CascadeMux
    port map (
            O => \N__4371\,
            I => \N__4368\
        );

    \I__963\ : InMux
    port map (
            O => \N__4368\,
            I => \N__4358\
        );

    \I__962\ : InMux
    port map (
            O => \N__4367\,
            I => \N__4343\
        );

    \I__961\ : InMux
    port map (
            O => \N__4366\,
            I => \N__4343\
        );

    \I__960\ : InMux
    port map (
            O => \N__4365\,
            I => \N__4343\
        );

    \I__959\ : InMux
    port map (
            O => \N__4364\,
            I => \N__4343\
        );

    \I__958\ : InMux
    port map (
            O => \N__4363\,
            I => \N__4343\
        );

    \I__957\ : InMux
    port map (
            O => \N__4362\,
            I => \N__4343\
        );

    \I__956\ : InMux
    port map (
            O => \N__4361\,
            I => \N__4343\
        );

    \I__955\ : LocalMux
    port map (
            O => \N__4358\,
            I => \N__4338\
        );

    \I__954\ : LocalMux
    port map (
            O => \N__4343\,
            I => \N__4335\
        );

    \I__953\ : InMux
    port map (
            O => \N__4342\,
            I => \N__4330\
        );

    \I__952\ : InMux
    port map (
            O => \N__4341\,
            I => \N__4330\
        );

    \I__951\ : Span4Mux_h
    port map (
            O => \N__4338\,
            I => \N__4323\
        );

    \I__950\ : Span4Mux_h
    port map (
            O => \N__4335\,
            I => \N__4323\
        );

    \I__949\ : LocalMux
    port map (
            O => \N__4330\,
            I => \N__4323\
        );

    \I__948\ : Odrv4
    port map (
            O => \N__4323\,
            I => n7_adj_1
        );

    \I__947\ : IoInMux
    port map (
            O => \N__4320\,
            I => \N__4317\
        );

    \I__946\ : LocalMux
    port map (
            O => \N__4317\,
            I => \N__4314\
        );

    \I__945\ : Span4Mux_s0_h
    port map (
            O => \N__4314\,
            I => \N__4310\
        );

    \I__944\ : InMux
    port map (
            O => \N__4313\,
            I => \N__4307\
        );

    \I__943\ : Span4Mux_v
    port map (
            O => \N__4310\,
            I => \N__4303\
        );

    \I__942\ : LocalMux
    port map (
            O => \N__4307\,
            I => \N__4300\
        );

    \I__941\ : InMux
    port map (
            O => \N__4306\,
            I => \N__4297\
        );

    \I__940\ : Odrv4
    port map (
            O => \N__4303\,
            I => io_leds_c_7
        );

    \I__939\ : Odrv12
    port map (
            O => \N__4300\,
            I => io_leds_c_7
        );

    \I__938\ : LocalMux
    port map (
            O => \N__4297\,
            I => io_leds_c_7
        );

    \I__937\ : InMux
    port map (
            O => \N__4290\,
            I => \N__4274\
        );

    \I__936\ : InMux
    port map (
            O => \N__4289\,
            I => \N__4274\
        );

    \I__935\ : InMux
    port map (
            O => \N__4288\,
            I => \N__4274\
        );

    \I__934\ : InMux
    port map (
            O => \N__4287\,
            I => \N__4274\
        );

    \I__933\ : InMux
    port map (
            O => \N__4286\,
            I => \N__4265\
        );

    \I__932\ : InMux
    port map (
            O => \N__4285\,
            I => \N__4265\
        );

    \I__931\ : InMux
    port map (
            O => \N__4284\,
            I => \N__4265\
        );

    \I__930\ : InMux
    port map (
            O => \N__4283\,
            I => \N__4265\
        );

    \I__929\ : LocalMux
    port map (
            O => \N__4274\,
            I => \N__4260\
        );

    \I__928\ : LocalMux
    port map (
            O => \N__4265\,
            I => \N__4260\
        );

    \I__927\ : Span4Mux_h
    port map (
            O => \N__4260\,
            I => \N__4257\
        );

    \I__926\ : Odrv4
    port map (
            O => \N__4257\,
            I => n7
        );

    \I__925\ : InMux
    port map (
            O => \N__4254\,
            I => \N__4250\
        );

    \I__924\ : CascadeMux
    port map (
            O => \N__4253\,
            I => \N__4247\
        );

    \I__923\ : LocalMux
    port map (
            O => \N__4250\,
            I => \N__4244\
        );

    \I__922\ : InMux
    port map (
            O => \N__4247\,
            I => \N__4241\
        );

    \I__921\ : Odrv4
    port map (
            O => \N__4244\,
            I => \ctrl_ledsArea_shifter_7\
        );

    \I__920\ : LocalMux
    port map (
            O => \N__4241\,
            I => \ctrl_ledsArea_shifter_7\
        );

    \I__919\ : CEMux
    port map (
            O => \N__4236\,
            I => \N__4233\
        );

    \I__918\ : LocalMux
    port map (
            O => \N__4233\,
            I => \N__4230\
        );

    \I__917\ : Span4Mux_h
    port map (
            O => \N__4230\,
            I => \N__4227\
        );

    \I__916\ : Odrv4
    port map (
            O => \N__4227\,
            I => n1353
        );

    \I__915\ : InMux
    port map (
            O => \N__4224\,
            I => \N__4210\
        );

    \I__914\ : InMux
    port map (
            O => \N__4223\,
            I => \N__4195\
        );

    \I__913\ : InMux
    port map (
            O => \N__4222\,
            I => \N__4195\
        );

    \I__912\ : InMux
    port map (
            O => \N__4221\,
            I => \N__4195\
        );

    \I__911\ : InMux
    port map (
            O => \N__4220\,
            I => \N__4195\
        );

    \I__910\ : InMux
    port map (
            O => \N__4219\,
            I => \N__4195\
        );

    \I__909\ : InMux
    port map (
            O => \N__4218\,
            I => \N__4195\
        );

    \I__908\ : InMux
    port map (
            O => \N__4217\,
            I => \N__4195\
        );

    \I__907\ : InMux
    port map (
            O => \N__4216\,
            I => \N__4192\
        );

    \I__906\ : InMux
    port map (
            O => \N__4215\,
            I => \N__4189\
        );

    \I__905\ : CascadeMux
    port map (
            O => \N__4214\,
            I => \N__4185\
        );

    \I__904\ : CascadeMux
    port map (
            O => \N__4213\,
            I => \N__4179\
        );

    \I__903\ : LocalMux
    port map (
            O => \N__4210\,
            I => \N__4161\
        );

    \I__902\ : LocalMux
    port map (
            O => \N__4195\,
            I => \N__4161\
        );

    \I__901\ : LocalMux
    port map (
            O => \N__4192\,
            I => \N__4161\
        );

    \I__900\ : LocalMux
    port map (
            O => \N__4189\,
            I => \N__4158\
        );

    \I__899\ : InMux
    port map (
            O => \N__4188\,
            I => \N__4151\
        );

    \I__898\ : InMux
    port map (
            O => \N__4185\,
            I => \N__4151\
        );

    \I__897\ : InMux
    port map (
            O => \N__4184\,
            I => \N__4151\
        );

    \I__896\ : InMux
    port map (
            O => \N__4183\,
            I => \N__4148\
        );

    \I__895\ : InMux
    port map (
            O => \N__4182\,
            I => \N__4141\
        );

    \I__894\ : InMux
    port map (
            O => \N__4179\,
            I => \N__4141\
        );

    \I__893\ : InMux
    port map (
            O => \N__4178\,
            I => \N__4138\
        );

    \I__892\ : InMux
    port map (
            O => \N__4177\,
            I => \N__4127\
        );

    \I__891\ : InMux
    port map (
            O => \N__4176\,
            I => \N__4127\
        );

    \I__890\ : InMux
    port map (
            O => \N__4175\,
            I => \N__4127\
        );

    \I__889\ : InMux
    port map (
            O => \N__4174\,
            I => \N__4127\
        );

    \I__888\ : InMux
    port map (
            O => \N__4173\,
            I => \N__4127\
        );

    \I__887\ : InMux
    port map (
            O => \N__4172\,
            I => \N__4116\
        );

    \I__886\ : InMux
    port map (
            O => \N__4171\,
            I => \N__4116\
        );

    \I__885\ : InMux
    port map (
            O => \N__4170\,
            I => \N__4116\
        );

    \I__884\ : InMux
    port map (
            O => \N__4169\,
            I => \N__4116\
        );

    \I__883\ : InMux
    port map (
            O => \N__4168\,
            I => \N__4116\
        );

    \I__882\ : Span4Mux_s3_v
    port map (
            O => \N__4161\,
            I => \N__4111\
        );

    \I__881\ : Span4Mux_v
    port map (
            O => \N__4158\,
            I => \N__4111\
        );

    \I__880\ : LocalMux
    port map (
            O => \N__4151\,
            I => \N__4106\
        );

    \I__879\ : LocalMux
    port map (
            O => \N__4148\,
            I => \N__4106\
        );

    \I__878\ : InMux
    port map (
            O => \N__4147\,
            I => \N__4101\
        );

    \I__877\ : InMux
    port map (
            O => \N__4146\,
            I => \N__4101\
        );

    \I__876\ : LocalMux
    port map (
            O => \N__4141\,
            I => ctrl_tap_fsm_state_0
        );

    \I__875\ : LocalMux
    port map (
            O => \N__4138\,
            I => ctrl_tap_fsm_state_0
        );

    \I__874\ : LocalMux
    port map (
            O => \N__4127\,
            I => ctrl_tap_fsm_state_0
        );

    \I__873\ : LocalMux
    port map (
            O => \N__4116\,
            I => ctrl_tap_fsm_state_0
        );

    \I__872\ : Odrv4
    port map (
            O => \N__4111\,
            I => ctrl_tap_fsm_state_0
        );

    \I__871\ : Odrv4
    port map (
            O => \N__4106\,
            I => ctrl_tap_fsm_state_0
        );

    \I__870\ : LocalMux
    port map (
            O => \N__4101\,
            I => ctrl_tap_fsm_state_0
        );

    \I__869\ : InMux
    port map (
            O => \N__4086\,
            I => \N__4080\
        );

    \I__868\ : InMux
    port map (
            O => \N__4085\,
            I => \N__4077\
        );

    \I__867\ : InMux
    port map (
            O => \N__4084\,
            I => \N__4073\
        );

    \I__866\ : CascadeMux
    port map (
            O => \N__4083\,
            I => \N__4059\
        );

    \I__865\ : LocalMux
    port map (
            O => \N__4080\,
            I => \N__4054\
        );

    \I__864\ : LocalMux
    port map (
            O => \N__4077\,
            I => \N__4054\
        );

    \I__863\ : InMux
    port map (
            O => \N__4076\,
            I => \N__4048\
        );

    \I__862\ : LocalMux
    port map (
            O => \N__4073\,
            I => \N__4045\
        );

    \I__861\ : InMux
    port map (
            O => \N__4072\,
            I => \N__4042\
        );

    \I__860\ : CascadeMux
    port map (
            O => \N__4071\,
            I => \N__4039\
        );

    \I__859\ : InMux
    port map (
            O => \N__4070\,
            I => \N__4033\
        );

    \I__858\ : InMux
    port map (
            O => \N__4069\,
            I => \N__4033\
        );

    \I__857\ : InMux
    port map (
            O => \N__4068\,
            I => \N__4030\
        );

    \I__856\ : InMux
    port map (
            O => \N__4067\,
            I => \N__4023\
        );

    \I__855\ : InMux
    port map (
            O => \N__4066\,
            I => \N__4023\
        );

    \I__854\ : InMux
    port map (
            O => \N__4065\,
            I => \N__4023\
        );

    \I__853\ : InMux
    port map (
            O => \N__4064\,
            I => \N__4014\
        );

    \I__852\ : InMux
    port map (
            O => \N__4063\,
            I => \N__4014\
        );

    \I__851\ : InMux
    port map (
            O => \N__4062\,
            I => \N__4014\
        );

    \I__850\ : InMux
    port map (
            O => \N__4059\,
            I => \N__4014\
        );

    \I__849\ : Span4Mux_h
    port map (
            O => \N__4054\,
            I => \N__4011\
        );

    \I__848\ : InMux
    port map (
            O => \N__4053\,
            I => \N__4004\
        );

    \I__847\ : InMux
    port map (
            O => \N__4052\,
            I => \N__4004\
        );

    \I__846\ : InMux
    port map (
            O => \N__4051\,
            I => \N__4004\
        );

    \I__845\ : LocalMux
    port map (
            O => \N__4048\,
            I => \N__3997\
        );

    \I__844\ : Span4Mux_h
    port map (
            O => \N__4045\,
            I => \N__3997\
        );

    \I__843\ : LocalMux
    port map (
            O => \N__4042\,
            I => \N__3997\
        );

    \I__842\ : InMux
    port map (
            O => \N__4039\,
            I => \N__3992\
        );

    \I__841\ : InMux
    port map (
            O => \N__4038\,
            I => \N__3992\
        );

    \I__840\ : LocalMux
    port map (
            O => \N__4033\,
            I => ctrl_tap_fsm_state_3
        );

    \I__839\ : LocalMux
    port map (
            O => \N__4030\,
            I => ctrl_tap_fsm_state_3
        );

    \I__838\ : LocalMux
    port map (
            O => \N__4023\,
            I => ctrl_tap_fsm_state_3
        );

    \I__837\ : LocalMux
    port map (
            O => \N__4014\,
            I => ctrl_tap_fsm_state_3
        );

    \I__836\ : Odrv4
    port map (
            O => \N__4011\,
            I => ctrl_tap_fsm_state_3
        );

    \I__835\ : LocalMux
    port map (
            O => \N__4004\,
            I => ctrl_tap_fsm_state_3
        );

    \I__834\ : Odrv4
    port map (
            O => \N__3997\,
            I => ctrl_tap_fsm_state_3
        );

    \I__833\ : LocalMux
    port map (
            O => \N__3992\,
            I => ctrl_tap_fsm_state_3
        );

    \I__832\ : CascadeMux
    port map (
            O => \N__3975\,
            I => \N__3969\
        );

    \I__831\ : CascadeMux
    port map (
            O => \N__3974\,
            I => \N__3965\
        );

    \I__830\ : CascadeMux
    port map (
            O => \N__3973\,
            I => \N__3958\
        );

    \I__829\ : InMux
    port map (
            O => \N__3972\,
            I => \N__3955\
        );

    \I__828\ : InMux
    port map (
            O => \N__3969\,
            I => \N__3950\
        );

    \I__827\ : InMux
    port map (
            O => \N__3968\,
            I => \N__3950\
        );

    \I__826\ : InMux
    port map (
            O => \N__3965\,
            I => \N__3945\
        );

    \I__825\ : InMux
    port map (
            O => \N__3964\,
            I => \N__3945\
        );

    \I__824\ : InMux
    port map (
            O => \N__3963\,
            I => \N__3938\
        );

    \I__823\ : InMux
    port map (
            O => \N__3962\,
            I => \N__3938\
        );

    \I__822\ : InMux
    port map (
            O => \N__3961\,
            I => \N__3938\
        );

    \I__821\ : InMux
    port map (
            O => \N__3958\,
            I => \N__3934\
        );

    \I__820\ : LocalMux
    port map (
            O => \N__3955\,
            I => \N__3930\
        );

    \I__819\ : LocalMux
    port map (
            O => \N__3950\,
            I => \N__3923\
        );

    \I__818\ : LocalMux
    port map (
            O => \N__3945\,
            I => \N__3923\
        );

    \I__817\ : LocalMux
    port map (
            O => \N__3938\,
            I => \N__3923\
        );

    \I__816\ : InMux
    port map (
            O => \N__3937\,
            I => \N__3920\
        );

    \I__815\ : LocalMux
    port map (
            O => \N__3934\,
            I => \N__3917\
        );

    \I__814\ : CascadeMux
    port map (
            O => \N__3933\,
            I => \N__3914\
        );

    \I__813\ : Span4Mux_v
    port map (
            O => \N__3930\,
            I => \N__3909\
        );

    \I__812\ : Span4Mux_v
    port map (
            O => \N__3923\,
            I => \N__3909\
        );

    \I__811\ : LocalMux
    port map (
            O => \N__3920\,
            I => \N__3906\
        );

    \I__810\ : Span4Mux_s3_h
    port map (
            O => \N__3917\,
            I => \N__3903\
        );

    \I__809\ : InMux
    port map (
            O => \N__3914\,
            I => \N__3900\
        );

    \I__808\ : IoSpan4Mux
    port map (
            O => \N__3909\,
            I => \N__3897\
        );

    \I__807\ : Span4Mux_s3_h
    port map (
            O => \N__3906\,
            I => \N__3894\
        );

    \I__806\ : Sp12to4
    port map (
            O => \N__3903\,
            I => \N__3889\
        );

    \I__805\ : LocalMux
    port map (
            O => \N__3900\,
            I => \N__3889\
        );

    \I__804\ : Odrv4
    port map (
            O => \N__3897\,
            I => \ctrl_tap_fsm_stateNext_3__N_10_c_3\
        );

    \I__803\ : Odrv4
    port map (
            O => \N__3894\,
            I => \ctrl_tap_fsm_stateNext_3__N_10_c_3\
        );

    \I__802\ : Odrv12
    port map (
            O => \N__3889\,
            I => \ctrl_tap_fsm_stateNext_3__N_10_c_3\
        );

    \I__801\ : InMux
    port map (
            O => \N__3882\,
            I => \N__3875\
        );

    \I__800\ : InMux
    port map (
            O => \N__3881\,
            I => \N__3875\
        );

    \I__799\ : InMux
    port map (
            O => \N__3880\,
            I => \N__3872\
        );

    \I__798\ : LocalMux
    port map (
            O => \N__3875\,
            I => \N__3865\
        );

    \I__797\ : LocalMux
    port map (
            O => \N__3872\,
            I => \N__3850\
        );

    \I__796\ : InMux
    port map (
            O => \N__3871\,
            I => \N__3843\
        );

    \I__795\ : InMux
    port map (
            O => \N__3870\,
            I => \N__3843\
        );

    \I__794\ : InMux
    port map (
            O => \N__3869\,
            I => \N__3843\
        );

    \I__793\ : InMux
    port map (
            O => \N__3868\,
            I => \N__3840\
        );

    \I__792\ : Span4Mux_h
    port map (
            O => \N__3865\,
            I => \N__3835\
        );

    \I__791\ : InMux
    port map (
            O => \N__3864\,
            I => \N__3832\
        );

    \I__790\ : InMux
    port map (
            O => \N__3863\,
            I => \N__3829\
        );

    \I__789\ : InMux
    port map (
            O => \N__3862\,
            I => \N__3818\
        );

    \I__788\ : InMux
    port map (
            O => \N__3861\,
            I => \N__3818\
        );

    \I__787\ : InMux
    port map (
            O => \N__3860\,
            I => \N__3818\
        );

    \I__786\ : InMux
    port map (
            O => \N__3859\,
            I => \N__3818\
        );

    \I__785\ : InMux
    port map (
            O => \N__3858\,
            I => \N__3818\
        );

    \I__784\ : InMux
    port map (
            O => \N__3857\,
            I => \N__3807\
        );

    \I__783\ : InMux
    port map (
            O => \N__3856\,
            I => \N__3807\
        );

    \I__782\ : InMux
    port map (
            O => \N__3855\,
            I => \N__3807\
        );

    \I__781\ : InMux
    port map (
            O => \N__3854\,
            I => \N__3807\
        );

    \I__780\ : InMux
    port map (
            O => \N__3853\,
            I => \N__3807\
        );

    \I__779\ : Span4Mux_h
    port map (
            O => \N__3850\,
            I => \N__3800\
        );

    \I__778\ : LocalMux
    port map (
            O => \N__3843\,
            I => \N__3800\
        );

    \I__777\ : LocalMux
    port map (
            O => \N__3840\,
            I => \N__3800\
        );

    \I__776\ : InMux
    port map (
            O => \N__3839\,
            I => \N__3795\
        );

    \I__775\ : InMux
    port map (
            O => \N__3838\,
            I => \N__3795\
        );

    \I__774\ : Odrv4
    port map (
            O => \N__3835\,
            I => ctrl_tap_fsm_state_1
        );

    \I__773\ : LocalMux
    port map (
            O => \N__3832\,
            I => ctrl_tap_fsm_state_1
        );

    \I__772\ : LocalMux
    port map (
            O => \N__3829\,
            I => ctrl_tap_fsm_state_1
        );

    \I__771\ : LocalMux
    port map (
            O => \N__3818\,
            I => ctrl_tap_fsm_state_1
        );

    \I__770\ : LocalMux
    port map (
            O => \N__3807\,
            I => ctrl_tap_fsm_state_1
        );

    \I__769\ : Odrv4
    port map (
            O => \N__3800\,
            I => ctrl_tap_fsm_state_1
        );

    \I__768\ : LocalMux
    port map (
            O => \N__3795\,
            I => ctrl_tap_fsm_state_1
        );

    \I__767\ : InMux
    port map (
            O => \N__3780\,
            I => \N__3777\
        );

    \I__766\ : LocalMux
    port map (
            O => \N__3777\,
            I => \N__3774\
        );

    \I__765\ : Span4Mux_s3_h
    port map (
            O => \N__3774\,
            I => \N__3771\
        );

    \I__764\ : Odrv4
    port map (
            O => \N__3771\,
            I => n963
        );

    \I__763\ : InMux
    port map (
            O => \N__3768\,
            I => \N__3765\
        );

    \I__762\ : LocalMux
    port map (
            O => \N__3765\,
            I => \N__3762\
        );

    \I__761\ : Span4Mux_h
    port map (
            O => \N__3762\,
            I => \N__3758\
        );

    \I__760\ : InMux
    port map (
            O => \N__3761\,
            I => \N__3755\
        );

    \I__759\ : Odrv4
    port map (
            O => \N__3758\,
            I => n15
        );

    \I__758\ : LocalMux
    port map (
            O => \N__3755\,
            I => n15
        );

    \I__757\ : CascadeMux
    port map (
            O => \N__3750\,
            I => \N__3747\
        );

    \I__756\ : InMux
    port map (
            O => \N__3747\,
            I => \N__3741\
        );

    \I__755\ : InMux
    port map (
            O => \N__3746\,
            I => \N__3741\
        );

    \I__754\ : LocalMux
    port map (
            O => \N__3741\,
            I => \ctrl_idcodeArea_shifter_18\
        );

    \I__753\ : CascadeMux
    port map (
            O => \N__3738\,
            I => \N__3734\
        );

    \I__752\ : InMux
    port map (
            O => \N__3737\,
            I => \N__3729\
        );

    \I__751\ : InMux
    port map (
            O => \N__3734\,
            I => \N__3729\
        );

    \I__750\ : LocalMux
    port map (
            O => \N__3729\,
            I => \ctrl_idcodeArea_shifter_20\
        );

    \I__749\ : InMux
    port map (
            O => \N__3726\,
            I => \N__3720\
        );

    \I__748\ : InMux
    port map (
            O => \N__3725\,
            I => \N__3720\
        );

    \I__747\ : LocalMux
    port map (
            O => \N__3720\,
            I => \ctrl_idcodeArea_shifter_19\
        );

    \I__746\ : InMux
    port map (
            O => \N__3717\,
            I => \N__3713\
        );

    \I__745\ : InMux
    port map (
            O => \N__3716\,
            I => \N__3710\
        );

    \I__744\ : LocalMux
    port map (
            O => \N__3713\,
            I => \N__3707\
        );

    \I__743\ : LocalMux
    port map (
            O => \N__3710\,
            I => \ctrl_idcodeArea_shifter_31\
        );

    \I__742\ : Odrv12
    port map (
            O => \N__3707\,
            I => \ctrl_idcodeArea_shifter_31\
        );

    \I__741\ : CascadeMux
    port map (
            O => \N__3702\,
            I => \N__3698\
        );

    \I__740\ : CascadeMux
    port map (
            O => \N__3701\,
            I => \N__3695\
        );

    \I__739\ : InMux
    port map (
            O => \N__3698\,
            I => \N__3685\
        );

    \I__738\ : InMux
    port map (
            O => \N__3695\,
            I => \N__3685\
        );

    \I__737\ : CascadeMux
    port map (
            O => \N__3694\,
            I => \N__3678\
        );

    \I__736\ : CascadeMux
    port map (
            O => \N__3693\,
            I => \N__3674\
        );

    \I__735\ : CascadeMux
    port map (
            O => \N__3692\,
            I => \N__3671\
        );

    \I__734\ : CascadeMux
    port map (
            O => \N__3691\,
            I => \N__3667\
        );

    \I__733\ : CascadeMux
    port map (
            O => \N__3690\,
            I => \N__3664\
        );

    \I__732\ : LocalMux
    port map (
            O => \N__3685\,
            I => \N__3660\
        );

    \I__731\ : InMux
    port map (
            O => \N__3684\,
            I => \N__3653\
        );

    \I__730\ : InMux
    port map (
            O => \N__3683\,
            I => \N__3653\
        );

    \I__729\ : InMux
    port map (
            O => \N__3682\,
            I => \N__3650\
        );

    \I__728\ : CascadeMux
    port map (
            O => \N__3681\,
            I => \N__3646\
        );

    \I__727\ : InMux
    port map (
            O => \N__3678\,
            I => \N__3641\
        );

    \I__726\ : InMux
    port map (
            O => \N__3677\,
            I => \N__3641\
        );

    \I__725\ : InMux
    port map (
            O => \N__3674\,
            I => \N__3636\
        );

    \I__724\ : InMux
    port map (
            O => \N__3671\,
            I => \N__3636\
        );

    \I__723\ : InMux
    port map (
            O => \N__3670\,
            I => \N__3627\
        );

    \I__722\ : InMux
    port map (
            O => \N__3667\,
            I => \N__3627\
        );

    \I__721\ : InMux
    port map (
            O => \N__3664\,
            I => \N__3627\
        );

    \I__720\ : InMux
    port map (
            O => \N__3663\,
            I => \N__3627\
        );

    \I__719\ : Span4Mux_h
    port map (
            O => \N__3660\,
            I => \N__3624\
        );

    \I__718\ : InMux
    port map (
            O => \N__3659\,
            I => \N__3619\
        );

    \I__717\ : InMux
    port map (
            O => \N__3658\,
            I => \N__3619\
        );

    \I__716\ : LocalMux
    port map (
            O => \N__3653\,
            I => \N__3614\
        );

    \I__715\ : LocalMux
    port map (
            O => \N__3650\,
            I => \N__3614\
        );

    \I__714\ : InMux
    port map (
            O => \N__3649\,
            I => \N__3609\
        );

    \I__713\ : InMux
    port map (
            O => \N__3646\,
            I => \N__3609\
        );

    \I__712\ : LocalMux
    port map (
            O => \N__3641\,
            I => ctrl_tap_fsm_state_2
        );

    \I__711\ : LocalMux
    port map (
            O => \N__3636\,
            I => ctrl_tap_fsm_state_2
        );

    \I__710\ : LocalMux
    port map (
            O => \N__3627\,
            I => ctrl_tap_fsm_state_2
        );

    \I__709\ : Odrv4
    port map (
            O => \N__3624\,
            I => ctrl_tap_fsm_state_2
        );

    \I__708\ : LocalMux
    port map (
            O => \N__3619\,
            I => ctrl_tap_fsm_state_2
        );

    \I__707\ : Odrv4
    port map (
            O => \N__3614\,
            I => ctrl_tap_fsm_state_2
        );

    \I__706\ : LocalMux
    port map (
            O => \N__3609\,
            I => ctrl_tap_fsm_state_2
        );

    \I__705\ : CEMux
    port map (
            O => \N__3594\,
            I => \N__3591\
        );

    \I__704\ : LocalMux
    port map (
            O => \N__3591\,
            I => \N__3587\
        );

    \I__703\ : CEMux
    port map (
            O => \N__3590\,
            I => \N__3584\
        );

    \I__702\ : Span4Mux_s1_v
    port map (
            O => \N__3587\,
            I => \N__3579\
        );

    \I__701\ : LocalMux
    port map (
            O => \N__3584\,
            I => \N__3579\
        );

    \I__700\ : Span4Mux_h
    port map (
            O => \N__3579\,
            I => \N__3576\
        );

    \I__699\ : Odrv4
    port map (
            O => \N__3576\,
            I => n1067
        );

    \I__698\ : CascadeMux
    port map (
            O => \N__3573\,
            I => \N__3570\
        );

    \I__697\ : InMux
    port map (
            O => \N__3570\,
            I => \N__3567\
        );

    \I__696\ : LocalMux
    port map (
            O => \N__3567\,
            I => \N__3563\
        );

    \I__695\ : InMux
    port map (
            O => \N__3566\,
            I => \N__3560\
        );

    \I__694\ : Odrv12
    port map (
            O => \N__3563\,
            I => \ctrl_idcodeArea_shifter_22\
        );

    \I__693\ : LocalMux
    port map (
            O => \N__3560\,
            I => \ctrl_idcodeArea_shifter_22\
        );

    \I__692\ : InMux
    port map (
            O => \N__3555\,
            I => \N__3549\
        );

    \I__691\ : InMux
    port map (
            O => \N__3554\,
            I => \N__3549\
        );

    \I__690\ : LocalMux
    port map (
            O => \N__3549\,
            I => \ctrl_idcodeArea_shifter_21\
        );

    \I__689\ : IoInMux
    port map (
            O => \N__3546\,
            I => \N__3543\
        );

    \I__688\ : LocalMux
    port map (
            O => \N__3543\,
            I => \N__3540\
        );

    \I__687\ : Span4Mux_s1_h
    port map (
            O => \N__3540\,
            I => \N__3536\
        );

    \I__686\ : InMux
    port map (
            O => \N__3539\,
            I => \N__3533\
        );

    \I__685\ : Sp12to4
    port map (
            O => \N__3536\,
            I => \N__3529\
        );

    \I__684\ : LocalMux
    port map (
            O => \N__3533\,
            I => \N__3526\
        );

    \I__683\ : InMux
    port map (
            O => \N__3532\,
            I => \N__3523\
        );

    \I__682\ : Span12Mux_v
    port map (
            O => \N__3529\,
            I => \N__3520\
        );

    \I__681\ : Span4Mux_v
    port map (
            O => \N__3526\,
            I => \N__3515\
        );

    \I__680\ : LocalMux
    port map (
            O => \N__3523\,
            I => \N__3515\
        );

    \I__679\ : Odrv12
    port map (
            O => \N__3520\,
            I => io_leds_c_0
        );

    \I__678\ : Odrv4
    port map (
            O => \N__3515\,
            I => io_leds_c_0
        );

    \I__677\ : InMux
    port map (
            O => \N__3510\,
            I => \N__3506\
        );

    \I__676\ : InMux
    port map (
            O => \N__3509\,
            I => \N__3503\
        );

    \I__675\ : LocalMux
    port map (
            O => \N__3506\,
            I => \N__3500\
        );

    \I__674\ : LocalMux
    port map (
            O => \N__3503\,
            I => \N__3497\
        );

    \I__673\ : Span4Mux_s3_v
    port map (
            O => \N__3500\,
            I => \N__3494\
        );

    \I__672\ : Span4Mux_s3_h
    port map (
            O => \N__3497\,
            I => \N__3491\
        );

    \I__671\ : Odrv4
    port map (
            O => \N__3494\,
            I => \ctrl_ledsArea_shifter_0\
        );

    \I__670\ : Odrv4
    port map (
            O => \N__3491\,
            I => \ctrl_ledsArea_shifter_0\
        );

    \I__669\ : SRMux
    port map (
            O => \N__3486\,
            I => \N__3482\
        );

    \I__668\ : SRMux
    port map (
            O => \N__3485\,
            I => \N__3479\
        );

    \I__667\ : LocalMux
    port map (
            O => \N__3482\,
            I => \N__3475\
        );

    \I__666\ : LocalMux
    port map (
            O => \N__3479\,
            I => \N__3472\
        );

    \I__665\ : SRMux
    port map (
            O => \N__3478\,
            I => \N__3469\
        );

    \I__664\ : Span4Mux_v
    port map (
            O => \N__3475\,
            I => \N__3464\
        );

    \I__663\ : Span4Mux_h
    port map (
            O => \N__3472\,
            I => \N__3464\
        );

    \I__662\ : LocalMux
    port map (
            O => \N__3469\,
            I => \N__3460\
        );

    \I__661\ : Span4Mux_v
    port map (
            O => \N__3464\,
            I => \N__3457\
        );

    \I__660\ : SRMux
    port map (
            O => \N__3463\,
            I => \N__3454\
        );

    \I__659\ : Span4Mux_v
    port map (
            O => \N__3460\,
            I => \N__3451\
        );

    \I__658\ : Span4Mux_v
    port map (
            O => \N__3457\,
            I => \N__3448\
        );

    \I__657\ : LocalMux
    port map (
            O => \N__3454\,
            I => \N__3445\
        );

    \I__656\ : Span4Mux_v
    port map (
            O => \N__3451\,
            I => \N__3442\
        );

    \I__655\ : Odrv4
    port map (
            O => \N__3448\,
            I => global_reset_c
        );

    \I__654\ : Odrv12
    port map (
            O => \N__3445\,
            I => global_reset_c
        );

    \I__653\ : Odrv4
    port map (
            O => \N__3442\,
            I => global_reset_c
        );

    \I__652\ : InMux
    port map (
            O => \N__3435\,
            I => \N__3432\
        );

    \I__651\ : LocalMux
    port map (
            O => \N__3432\,
            I => \N__3425\
        );

    \I__650\ : InMux
    port map (
            O => \N__3431\,
            I => \N__3422\
        );

    \I__649\ : InMux
    port map (
            O => \N__3430\,
            I => \N__3417\
        );

    \I__648\ : InMux
    port map (
            O => \N__3429\,
            I => \N__3417\
        );

    \I__647\ : InMux
    port map (
            O => \N__3428\,
            I => \N__3414\
        );

    \I__646\ : Odrv4
    port map (
            O => \N__3425\,
            I => ctrl_tap_instruction_1
        );

    \I__645\ : LocalMux
    port map (
            O => \N__3422\,
            I => ctrl_tap_instruction_1
        );

    \I__644\ : LocalMux
    port map (
            O => \N__3417\,
            I => ctrl_tap_instruction_1
        );

    \I__643\ : LocalMux
    port map (
            O => \N__3414\,
            I => ctrl_tap_instruction_1
        );

    \I__642\ : CascadeMux
    port map (
            O => \N__3405\,
            I => \N__3401\
        );

    \I__641\ : InMux
    port map (
            O => \N__3404\,
            I => \N__3398\
        );

    \I__640\ : InMux
    port map (
            O => \N__3401\,
            I => \N__3393\
        );

    \I__639\ : LocalMux
    port map (
            O => \N__3398\,
            I => \N__3390\
        );

    \I__638\ : InMux
    port map (
            O => \N__3397\,
            I => \N__3387\
        );

    \I__637\ : InMux
    port map (
            O => \N__3396\,
            I => \N__3384\
        );

    \I__636\ : LocalMux
    port map (
            O => \N__3393\,
            I => ctrl_tap_instruction_2
        );

    \I__635\ : Odrv4
    port map (
            O => \N__3390\,
            I => ctrl_tap_instruction_2
        );

    \I__634\ : LocalMux
    port map (
            O => \N__3387\,
            I => ctrl_tap_instruction_2
        );

    \I__633\ : LocalMux
    port map (
            O => \N__3384\,
            I => ctrl_tap_instruction_2
        );

    \I__632\ : InMux
    port map (
            O => \N__3375\,
            I => \N__3372\
        );

    \I__631\ : LocalMux
    port map (
            O => \N__3372\,
            I => \N__3368\
        );

    \I__630\ : InMux
    port map (
            O => \N__3371\,
            I => \N__3365\
        );

    \I__629\ : Odrv12
    port map (
            O => \N__3368\,
            I => \ctrl_tap_instructionShift_2\
        );

    \I__628\ : LocalMux
    port map (
            O => \N__3365\,
            I => \ctrl_tap_instructionShift_2\
        );

    \I__627\ : InMux
    port map (
            O => \N__3360\,
            I => \N__3356\
        );

    \I__626\ : InMux
    port map (
            O => \N__3359\,
            I => \N__3353\
        );

    \I__625\ : LocalMux
    port map (
            O => \N__3356\,
            I => \N__3347\
        );

    \I__624\ : LocalMux
    port map (
            O => \N__3353\,
            I => \N__3347\
        );

    \I__623\ : InMux
    port map (
            O => \N__3352\,
            I => \N__3344\
        );

    \I__622\ : Odrv4
    port map (
            O => \N__3347\,
            I => ctrl_tap_instruction_4
        );

    \I__621\ : LocalMux
    port map (
            O => \N__3344\,
            I => ctrl_tap_instruction_4
        );

    \I__620\ : InMux
    port map (
            O => \N__3339\,
            I => \N__3336\
        );

    \I__619\ : LocalMux
    port map (
            O => \N__3336\,
            I => \N__3331\
        );

    \I__618\ : InMux
    port map (
            O => \N__3335\,
            I => \N__3326\
        );

    \I__617\ : InMux
    port map (
            O => \N__3334\,
            I => \N__3326\
        );

    \I__616\ : Odrv12
    port map (
            O => \N__3331\,
            I => ctrl_tap_instruction_5
        );

    \I__615\ : LocalMux
    port map (
            O => \N__3326\,
            I => ctrl_tap_instruction_5
        );

    \I__614\ : CascadeMux
    port map (
            O => \N__3321\,
            I => \N__3318\
        );

    \I__613\ : InMux
    port map (
            O => \N__3318\,
            I => \N__3315\
        );

    \I__612\ : LocalMux
    port map (
            O => \N__3315\,
            I => \N__3312\
        );

    \I__611\ : Span4Mux_s2_h
    port map (
            O => \N__3312\,
            I => \N__3308\
        );

    \I__610\ : InMux
    port map (
            O => \N__3311\,
            I => \N__3305\
        );

    \I__609\ : Odrv4
    port map (
            O => \N__3308\,
            I => \ctrl_tap_instructionShift_5\
        );

    \I__608\ : LocalMux
    port map (
            O => \N__3305\,
            I => \ctrl_tap_instructionShift_5\
        );

    \I__607\ : CascadeMux
    port map (
            O => \N__3300\,
            I => \N__3296\
        );

    \I__606\ : InMux
    port map (
            O => \N__3299\,
            I => \N__3293\
        );

    \I__605\ : InMux
    port map (
            O => \N__3296\,
            I => \N__3288\
        );

    \I__604\ : LocalMux
    port map (
            O => \N__3293\,
            I => \N__3285\
        );

    \I__603\ : InMux
    port map (
            O => \N__3292\,
            I => \N__3280\
        );

    \I__602\ : InMux
    port map (
            O => \N__3291\,
            I => \N__3280\
        );

    \I__601\ : LocalMux
    port map (
            O => \N__3288\,
            I => ctrl_tap_instruction_7
        );

    \I__600\ : Odrv4
    port map (
            O => \N__3285\,
            I => ctrl_tap_instruction_7
        );

    \I__599\ : LocalMux
    port map (
            O => \N__3280\,
            I => ctrl_tap_instruction_7
        );

    \I__598\ : CascadeMux
    port map (
            O => \N__3273\,
            I => \N__3270\
        );

    \I__597\ : InMux
    port map (
            O => \N__3270\,
            I => \N__3267\
        );

    \I__596\ : LocalMux
    port map (
            O => \N__3267\,
            I => \N__3264\
        );

    \I__595\ : Span4Mux_s2_h
    port map (
            O => \N__3264\,
            I => \N__3260\
        );

    \I__594\ : InMux
    port map (
            O => \N__3263\,
            I => \N__3257\
        );

    \I__593\ : Odrv4
    port map (
            O => \N__3260\,
            I => \ctrl_tap_instructionShift_4\
        );

    \I__592\ : LocalMux
    port map (
            O => \N__3257\,
            I => \ctrl_tap_instructionShift_4\
        );

    \I__591\ : InMux
    port map (
            O => \N__3252\,
            I => \N__3248\
        );

    \I__590\ : CascadeMux
    port map (
            O => \N__3251\,
            I => \N__3244\
        );

    \I__589\ : LocalMux
    port map (
            O => \N__3248\,
            I => \N__3240\
        );

    \I__588\ : InMux
    port map (
            O => \N__3247\,
            I => \N__3237\
        );

    \I__587\ : InMux
    port map (
            O => \N__3244\,
            I => \N__3232\
        );

    \I__586\ : InMux
    port map (
            O => \N__3243\,
            I => \N__3232\
        );

    \I__585\ : Odrv4
    port map (
            O => \N__3240\,
            I => ctrl_tap_instruction_3
        );

    \I__584\ : LocalMux
    port map (
            O => \N__3237\,
            I => ctrl_tap_instruction_3
        );

    \I__583\ : LocalMux
    port map (
            O => \N__3232\,
            I => ctrl_tap_instruction_3
        );

    \I__582\ : CascadeMux
    port map (
            O => \N__3225\,
            I => \N__3222\
        );

    \I__581\ : InMux
    port map (
            O => \N__3222\,
            I => \N__3219\
        );

    \I__580\ : LocalMux
    port map (
            O => \N__3219\,
            I => \N__3215\
        );

    \I__579\ : InMux
    port map (
            O => \N__3218\,
            I => \N__3212\
        );

    \I__578\ : Odrv4
    port map (
            O => \N__3215\,
            I => \ctrl_tap_instructionShift_3\
        );

    \I__577\ : LocalMux
    port map (
            O => \N__3212\,
            I => \ctrl_tap_instructionShift_3\
        );

    \I__576\ : InMux
    port map (
            O => \N__3207\,
            I => \N__3204\
        );

    \I__575\ : LocalMux
    port map (
            O => \N__3204\,
            I => \N__3200\
        );

    \I__574\ : InMux
    port map (
            O => \N__3203\,
            I => \N__3197\
        );

    \I__573\ : Odrv4
    port map (
            O => \N__3200\,
            I => \ctrl_tap_instructionShift_7\
        );

    \I__572\ : LocalMux
    port map (
            O => \N__3197\,
            I => \ctrl_tap_instructionShift_7\
        );

    \I__571\ : InMux
    port map (
            O => \N__3192\,
            I => \N__3189\
        );

    \I__570\ : LocalMux
    port map (
            O => \N__3189\,
            I => \N__3183\
        );

    \I__569\ : InMux
    port map (
            O => \N__3188\,
            I => \N__3176\
        );

    \I__568\ : InMux
    port map (
            O => \N__3187\,
            I => \N__3176\
        );

    \I__567\ : InMux
    port map (
            O => \N__3186\,
            I => \N__3176\
        );

    \I__566\ : Odrv12
    port map (
            O => \N__3183\,
            I => ctrl_tap_instruction_6
        );

    \I__565\ : LocalMux
    port map (
            O => \N__3176\,
            I => ctrl_tap_instruction_6
        );

    \I__564\ : CascadeMux
    port map (
            O => \N__3171\,
            I => \N__3168\
        );

    \I__563\ : InMux
    port map (
            O => \N__3168\,
            I => \N__3165\
        );

    \I__562\ : LocalMux
    port map (
            O => \N__3165\,
            I => \N__3161\
        );

    \I__561\ : InMux
    port map (
            O => \N__3164\,
            I => \N__3158\
        );

    \I__560\ : Odrv4
    port map (
            O => \N__3161\,
            I => \ctrl_tap_instructionShift_6\
        );

    \I__559\ : LocalMux
    port map (
            O => \N__3158\,
            I => \ctrl_tap_instructionShift_6\
        );

    \I__558\ : CascadeMux
    port map (
            O => \N__3153\,
            I => \N__3150\
        );

    \I__557\ : InMux
    port map (
            O => \N__3150\,
            I => \N__3147\
        );

    \I__556\ : LocalMux
    port map (
            O => \N__3147\,
            I => \N__3143\
        );

    \I__555\ : InMux
    port map (
            O => \N__3146\,
            I => \N__3140\
        );

    \I__554\ : Odrv12
    port map (
            O => \N__3143\,
            I => \ctrl_tap_instructionShift_1\
        );

    \I__553\ : LocalMux
    port map (
            O => \N__3140\,
            I => \ctrl_tap_instructionShift_1\
        );

    \I__552\ : InMux
    port map (
            O => \N__3135\,
            I => \N__3132\
        );

    \I__551\ : LocalMux
    port map (
            O => \N__3132\,
            I => \N__3129\
        );

    \I__550\ : Span4Mux_h
    port map (
            O => \N__3129\,
            I => \N__3122\
        );

    \I__549\ : InMux
    port map (
            O => \N__3128\,
            I => \N__3119\
        );

    \I__548\ : InMux
    port map (
            O => \N__3127\,
            I => \N__3116\
        );

    \I__547\ : InMux
    port map (
            O => \N__3126\,
            I => \N__3113\
        );

    \I__546\ : InMux
    port map (
            O => \N__3125\,
            I => \N__3110\
        );

    \I__545\ : Odrv4
    port map (
            O => \N__3122\,
            I => ctrl_tap_instruction_0
        );

    \I__544\ : LocalMux
    port map (
            O => \N__3119\,
            I => ctrl_tap_instruction_0
        );

    \I__543\ : LocalMux
    port map (
            O => \N__3116\,
            I => ctrl_tap_instruction_0
        );

    \I__542\ : LocalMux
    port map (
            O => \N__3113\,
            I => ctrl_tap_instruction_0
        );

    \I__541\ : LocalMux
    port map (
            O => \N__3110\,
            I => ctrl_tap_instruction_0
        );

    \I__540\ : CascadeMux
    port map (
            O => \N__3099\,
            I => \N__3096\
        );

    \I__539\ : InMux
    port map (
            O => \N__3096\,
            I => \N__3093\
        );

    \I__538\ : LocalMux
    port map (
            O => \N__3093\,
            I => \N__3089\
        );

    \I__537\ : InMux
    port map (
            O => \N__3092\,
            I => \N__3086\
        );

    \I__536\ : Span4Mux_s1_v
    port map (
            O => \N__3089\,
            I => \N__3081\
        );

    \I__535\ : LocalMux
    port map (
            O => \N__3086\,
            I => \N__3081\
        );

    \I__534\ : Odrv4
    port map (
            O => \N__3081\,
            I => \ctrl_tap_instructionShift_0\
        );

    \I__533\ : CascadeMux
    port map (
            O => \N__3078\,
            I => \N__3075\
        );

    \I__532\ : InMux
    port map (
            O => \N__3075\,
            I => \N__3069\
        );

    \I__531\ : InMux
    port map (
            O => \N__3074\,
            I => \N__3069\
        );

    \I__530\ : LocalMux
    port map (
            O => \N__3069\,
            I => \ctrl_idcodeArea_shifter_11\
        );

    \I__529\ : InMux
    port map (
            O => \N__3066\,
            I => \N__3060\
        );

    \I__528\ : InMux
    port map (
            O => \N__3065\,
            I => \N__3060\
        );

    \I__527\ : LocalMux
    port map (
            O => \N__3060\,
            I => \ctrl_idcodeArea_shifter_10\
        );

    \I__526\ : InMux
    port map (
            O => \N__3057\,
            I => \N__3053\
        );

    \I__525\ : InMux
    port map (
            O => \N__3056\,
            I => \N__3050\
        );

    \I__524\ : LocalMux
    port map (
            O => \N__3053\,
            I => \myClockArea_timeout_counter_value_4\
        );

    \I__523\ : LocalMux
    port map (
            O => \N__3050\,
            I => \myClockArea_timeout_counter_value_4\
        );

    \I__522\ : InMux
    port map (
            O => \N__3045\,
            I => \N__3041\
        );

    \I__521\ : InMux
    port map (
            O => \N__3044\,
            I => \N__3038\
        );

    \I__520\ : LocalMux
    port map (
            O => \N__3041\,
            I => \myClockArea_timeout_counter_value_6\
        );

    \I__519\ : LocalMux
    port map (
            O => \N__3038\,
            I => \myClockArea_timeout_counter_value_6\
        );

    \I__518\ : CascadeMux
    port map (
            O => \N__3033\,
            I => \N__3029\
        );

    \I__517\ : InMux
    port map (
            O => \N__3032\,
            I => \N__3026\
        );

    \I__516\ : InMux
    port map (
            O => \N__3029\,
            I => \N__3023\
        );

    \I__515\ : LocalMux
    port map (
            O => \N__3026\,
            I => \myClockArea_timeout_counter_value_22\
        );

    \I__514\ : LocalMux
    port map (
            O => \N__3023\,
            I => \myClockArea_timeout_counter_value_22\
        );

    \I__513\ : InMux
    port map (
            O => \N__3018\,
            I => \N__3014\
        );

    \I__512\ : InMux
    port map (
            O => \N__3017\,
            I => \N__3011\
        );

    \I__511\ : LocalMux
    port map (
            O => \N__3014\,
            I => \myClockArea_timeout_counter_value_16\
        );

    \I__510\ : LocalMux
    port map (
            O => \N__3011\,
            I => \myClockArea_timeout_counter_value_16\
        );

    \I__509\ : InMux
    port map (
            O => \N__3006\,
            I => \N__3002\
        );

    \I__508\ : InMux
    port map (
            O => \N__3005\,
            I => \N__2999\
        );

    \I__507\ : LocalMux
    port map (
            O => \N__3002\,
            I => \myClockArea_timeout_counter_value_17\
        );

    \I__506\ : LocalMux
    port map (
            O => \N__2999\,
            I => \myClockArea_timeout_counter_value_17\
        );

    \I__505\ : InMux
    port map (
            O => \N__2994\,
            I => \N__2990\
        );

    \I__504\ : InMux
    port map (
            O => \N__2993\,
            I => \N__2987\
        );

    \I__503\ : LocalMux
    port map (
            O => \N__2990\,
            I => \myClockArea_timeout_counter_value_8\
        );

    \I__502\ : LocalMux
    port map (
            O => \N__2987\,
            I => \myClockArea_timeout_counter_value_8\
        );

    \I__501\ : CascadeMux
    port map (
            O => \N__2982\,
            I => \N__2978\
        );

    \I__500\ : InMux
    port map (
            O => \N__2981\,
            I => \N__2975\
        );

    \I__499\ : InMux
    port map (
            O => \N__2978\,
            I => \N__2972\
        );

    \I__498\ : LocalMux
    port map (
            O => \N__2975\,
            I => \myClockArea_timeout_counter_value_10\
        );

    \I__497\ : LocalMux
    port map (
            O => \N__2972\,
            I => \myClockArea_timeout_counter_value_10\
        );

    \I__496\ : InMux
    port map (
            O => \N__2967\,
            I => \N__2963\
        );

    \I__495\ : InMux
    port map (
            O => \N__2966\,
            I => \N__2960\
        );

    \I__494\ : LocalMux
    port map (
            O => \N__2963\,
            I => \myClockArea_timeout_counter_value_2\
        );

    \I__493\ : LocalMux
    port map (
            O => \N__2960\,
            I => \myClockArea_timeout_counter_value_2\
        );

    \I__492\ : InMux
    port map (
            O => \N__2955\,
            I => \N__2952\
        );

    \I__491\ : LocalMux
    port map (
            O => \N__2952\,
            I => n2176
        );

    \I__490\ : CascadeMux
    port map (
            O => \N__2949\,
            I => \n2160_cascade_\
        );

    \I__489\ : InMux
    port map (
            O => \N__2946\,
            I => \N__2943\
        );

    \I__488\ : LocalMux
    port map (
            O => \N__2943\,
            I => n2164
        );

    \I__487\ : InMux
    port map (
            O => \N__2940\,
            I => \N__2936\
        );

    \I__486\ : InMux
    port map (
            O => \N__2939\,
            I => \N__2933\
        );

    \I__485\ : LocalMux
    port map (
            O => \N__2936\,
            I => \myClockArea_timeout_counter_value_13\
        );

    \I__484\ : LocalMux
    port map (
            O => \N__2933\,
            I => \myClockArea_timeout_counter_value_13\
        );

    \I__483\ : InMux
    port map (
            O => \N__2928\,
            I => \N__2925\
        );

    \I__482\ : LocalMux
    port map (
            O => \N__2925\,
            I => n11
        );

    \I__481\ : CascadeMux
    port map (
            O => \N__2922\,
            I => \n2182_cascade_\
        );

    \I__480\ : InMux
    port map (
            O => \N__2919\,
            I => \N__2916\
        );

    \I__479\ : LocalMux
    port map (
            O => \N__2916\,
            I => n13
        );

    \I__478\ : CascadeMux
    port map (
            O => \N__2913\,
            I => \n2113_cascade_\
        );

    \I__477\ : InMux
    port map (
            O => \N__2910\,
            I => \N__2890\
        );

    \I__476\ : InMux
    port map (
            O => \N__2909\,
            I => \N__2890\
        );

    \I__475\ : InMux
    port map (
            O => \N__2908\,
            I => \N__2890\
        );

    \I__474\ : InMux
    port map (
            O => \N__2907\,
            I => \N__2890\
        );

    \I__473\ : InMux
    port map (
            O => \N__2906\,
            I => \N__2881\
        );

    \I__472\ : InMux
    port map (
            O => \N__2905\,
            I => \N__2881\
        );

    \I__471\ : InMux
    port map (
            O => \N__2904\,
            I => \N__2881\
        );

    \I__470\ : InMux
    port map (
            O => \N__2903\,
            I => \N__2881\
        );

    \I__469\ : InMux
    port map (
            O => \N__2902\,
            I => \N__2861\
        );

    \I__468\ : InMux
    port map (
            O => \N__2901\,
            I => \N__2861\
        );

    \I__467\ : InMux
    port map (
            O => \N__2900\,
            I => \N__2861\
        );

    \I__466\ : InMux
    port map (
            O => \N__2899\,
            I => \N__2861\
        );

    \I__465\ : LocalMux
    port map (
            O => \N__2890\,
            I => \N__2858\
        );

    \I__464\ : LocalMux
    port map (
            O => \N__2881\,
            I => \N__2855\
        );

    \I__463\ : InMux
    port map (
            O => \N__2880\,
            I => \N__2846\
        );

    \I__462\ : InMux
    port map (
            O => \N__2879\,
            I => \N__2846\
        );

    \I__461\ : InMux
    port map (
            O => \N__2878\,
            I => \N__2846\
        );

    \I__460\ : InMux
    port map (
            O => \N__2877\,
            I => \N__2846\
        );

    \I__459\ : InMux
    port map (
            O => \N__2876\,
            I => \N__2839\
        );

    \I__458\ : InMux
    port map (
            O => \N__2875\,
            I => \N__2839\
        );

    \I__457\ : InMux
    port map (
            O => \N__2874\,
            I => \N__2839\
        );

    \I__456\ : InMux
    port map (
            O => \N__2873\,
            I => \N__2830\
        );

    \I__455\ : InMux
    port map (
            O => \N__2872\,
            I => \N__2830\
        );

    \I__454\ : InMux
    port map (
            O => \N__2871\,
            I => \N__2830\
        );

    \I__453\ : InMux
    port map (
            O => \N__2870\,
            I => \N__2830\
        );

    \I__452\ : LocalMux
    port map (
            O => \N__2861\,
            I => n1771
        );

    \I__451\ : Odrv4
    port map (
            O => \N__2858\,
            I => n1771
        );

    \I__450\ : Odrv4
    port map (
            O => \N__2855\,
            I => n1771
        );

    \I__449\ : LocalMux
    port map (
            O => \N__2846\,
            I => n1771
        );

    \I__448\ : LocalMux
    port map (
            O => \N__2839\,
            I => n1771
        );

    \I__447\ : LocalMux
    port map (
            O => \N__2830\,
            I => n1771
        );

    \I__446\ : InMux
    port map (
            O => \N__2817\,
            I => \N__2813\
        );

    \I__445\ : InMux
    port map (
            O => \N__2816\,
            I => \N__2810\
        );

    \I__444\ : LocalMux
    port map (
            O => \N__2813\,
            I => \myClockArea_timeout_counter_value_19\
        );

    \I__443\ : LocalMux
    port map (
            O => \N__2810\,
            I => \myClockArea_timeout_counter_value_19\
        );

    \I__442\ : InMux
    port map (
            O => \N__2805\,
            I => \N__2801\
        );

    \I__441\ : InMux
    port map (
            O => \N__2804\,
            I => \N__2798\
        );

    \I__440\ : LocalMux
    port map (
            O => \N__2801\,
            I => \myClockArea_timeout_counter_value_15\
        );

    \I__439\ : LocalMux
    port map (
            O => \N__2798\,
            I => \myClockArea_timeout_counter_value_15\
        );

    \I__438\ : CascadeMux
    port map (
            O => \N__2793\,
            I => \N__2789\
        );

    \I__437\ : InMux
    port map (
            O => \N__2792\,
            I => \N__2786\
        );

    \I__436\ : InMux
    port map (
            O => \N__2789\,
            I => \N__2783\
        );

    \I__435\ : LocalMux
    port map (
            O => \N__2786\,
            I => \myClockArea_timeout_counter_value_20\
        );

    \I__434\ : LocalMux
    port map (
            O => \N__2783\,
            I => \myClockArea_timeout_counter_value_20\
        );

    \I__433\ : InMux
    port map (
            O => \N__2778\,
            I => \N__2774\
        );

    \I__432\ : InMux
    port map (
            O => \N__2777\,
            I => \N__2771\
        );

    \I__431\ : LocalMux
    port map (
            O => \N__2774\,
            I => \myClockArea_timeout_counter_value_11\
        );

    \I__430\ : LocalMux
    port map (
            O => \N__2771\,
            I => \myClockArea_timeout_counter_value_11\
        );

    \I__429\ : InMux
    port map (
            O => \N__2766\,
            I => \N__2763\
        );

    \I__428\ : LocalMux
    port map (
            O => \N__2763\,
            I => n2162
        );

    \I__427\ : InMux
    port map (
            O => \N__2760\,
            I => \N__2757\
        );

    \I__426\ : LocalMux
    port map (
            O => \N__2757\,
            I => n2113
        );

    \I__425\ : InMux
    port map (
            O => \N__2754\,
            I => \N__2737\
        );

    \I__424\ : InMux
    port map (
            O => \N__2753\,
            I => \N__2737\
        );

    \I__423\ : InMux
    port map (
            O => \N__2752\,
            I => \N__2737\
        );

    \I__422\ : InMux
    port map (
            O => \N__2751\,
            I => \N__2737\
        );

    \I__421\ : InMux
    port map (
            O => \N__2750\,
            I => \N__2737\
        );

    \I__420\ : InMux
    port map (
            O => \N__2749\,
            I => \N__2734\
        );

    \I__419\ : InMux
    port map (
            O => \N__2748\,
            I => \N__2731\
        );

    \I__418\ : LocalMux
    port map (
            O => \N__2737\,
            I => n12_adj_3
        );

    \I__417\ : LocalMux
    port map (
            O => \N__2734\,
            I => n12_adj_3
        );

    \I__416\ : LocalMux
    port map (
            O => \N__2731\,
            I => n12_adj_3
        );

    \I__415\ : InMux
    port map (
            O => \N__2724\,
            I => \N__2712\
        );

    \I__414\ : InMux
    port map (
            O => \N__2723\,
            I => \N__2712\
        );

    \I__413\ : InMux
    port map (
            O => \N__2722\,
            I => \N__2712\
        );

    \I__412\ : InMux
    port map (
            O => \N__2721\,
            I => \N__2712\
        );

    \I__411\ : LocalMux
    port map (
            O => \N__2712\,
            I => n1769
        );

    \I__410\ : InMux
    port map (
            O => \N__2709\,
            I => \N__2706\
        );

    \I__409\ : LocalMux
    port map (
            O => \N__2706\,
            I => n1864
        );

    \I__408\ : InMux
    port map (
            O => \N__2703\,
            I => \N__2699\
        );

    \I__407\ : InMux
    port map (
            O => \N__2702\,
            I => \N__2696\
        );

    \I__406\ : LocalMux
    port map (
            O => \N__2699\,
            I => \myClockArea_timeout_counter_value_3\
        );

    \I__405\ : LocalMux
    port map (
            O => \N__2696\,
            I => \myClockArea_timeout_counter_value_3\
        );

    \I__404\ : InMux
    port map (
            O => \N__2691\,
            I => \N__2687\
        );

    \I__403\ : InMux
    port map (
            O => \N__2690\,
            I => \N__2684\
        );

    \I__402\ : LocalMux
    port map (
            O => \N__2687\,
            I => \myClockArea_timeout_counter_value_1\
        );

    \I__401\ : LocalMux
    port map (
            O => \N__2684\,
            I => \myClockArea_timeout_counter_value_1\
        );

    \I__400\ : CascadeMux
    port map (
            O => \N__2679\,
            I => \N__2675\
        );

    \I__399\ : InMux
    port map (
            O => \N__2678\,
            I => \N__2672\
        );

    \I__398\ : InMux
    port map (
            O => \N__2675\,
            I => \N__2669\
        );

    \I__397\ : LocalMux
    port map (
            O => \N__2672\,
            I => \myClockArea_timeout_counter_value_5\
        );

    \I__396\ : LocalMux
    port map (
            O => \N__2669\,
            I => \myClockArea_timeout_counter_value_5\
        );

    \I__395\ : InMux
    port map (
            O => \N__2664\,
            I => \N__2660\
        );

    \I__394\ : InMux
    port map (
            O => \N__2663\,
            I => \N__2657\
        );

    \I__393\ : LocalMux
    port map (
            O => \N__2660\,
            I => \myClockArea_timeout_counter_value_0\
        );

    \I__392\ : LocalMux
    port map (
            O => \N__2657\,
            I => \myClockArea_timeout_counter_value_0\
        );

    \I__391\ : InMux
    port map (
            O => \N__2652\,
            I => \N__2648\
        );

    \I__390\ : InMux
    port map (
            O => \N__2651\,
            I => \N__2645\
        );

    \I__389\ : LocalMux
    port map (
            O => \N__2648\,
            I => \myClockArea_timeout_counter_value_9\
        );

    \I__388\ : LocalMux
    port map (
            O => \N__2645\,
            I => \myClockArea_timeout_counter_value_9\
        );

    \I__387\ : InMux
    port map (
            O => \N__2640\,
            I => \N__2636\
        );

    \I__386\ : InMux
    port map (
            O => \N__2639\,
            I => \N__2633\
        );

    \I__385\ : LocalMux
    port map (
            O => \N__2636\,
            I => \N__2630\
        );

    \I__384\ : LocalMux
    port map (
            O => \N__2633\,
            I => \myClockArea_timeout_counter_value_18\
        );

    \I__383\ : Odrv4
    port map (
            O => \N__2630\,
            I => \myClockArea_timeout_counter_value_18\
        );

    \I__382\ : CascadeMux
    port map (
            O => \N__2625\,
            I => \N__2621\
        );

    \I__381\ : InMux
    port map (
            O => \N__2624\,
            I => \N__2618\
        );

    \I__380\ : InMux
    port map (
            O => \N__2621\,
            I => \N__2615\
        );

    \I__379\ : LocalMux
    port map (
            O => \N__2618\,
            I => \myClockArea_timeout_counter_value_12\
        );

    \I__378\ : LocalMux
    port map (
            O => \N__2615\,
            I => \myClockArea_timeout_counter_value_12\
        );

    \I__377\ : InMux
    port map (
            O => \N__2610\,
            I => \N__2606\
        );

    \I__376\ : InMux
    port map (
            O => \N__2609\,
            I => \N__2603\
        );

    \I__375\ : LocalMux
    port map (
            O => \N__2606\,
            I => \myClockArea_timeout_counter_value_14\
        );

    \I__374\ : LocalMux
    port map (
            O => \N__2603\,
            I => \myClockArea_timeout_counter_value_14\
        );

    \I__373\ : CascadeMux
    port map (
            O => \N__2598\,
            I => \N__2594\
        );

    \I__372\ : InMux
    port map (
            O => \N__2597\,
            I => \N__2591\
        );

    \I__371\ : InMux
    port map (
            O => \N__2594\,
            I => \N__2588\
        );

    \I__370\ : LocalMux
    port map (
            O => \N__2591\,
            I => \ctrl_idcodeArea_shifter_9\
        );

    \I__369\ : LocalMux
    port map (
            O => \N__2588\,
            I => \ctrl_idcodeArea_shifter_9\
        );

    \I__368\ : InMux
    port map (
            O => \N__2583\,
            I => \N__2579\
        );

    \I__367\ : InMux
    port map (
            O => \N__2582\,
            I => \N__2576\
        );

    \I__366\ : LocalMux
    port map (
            O => \N__2579\,
            I => \myClockArea_timeout_counter_value_7\
        );

    \I__365\ : LocalMux
    port map (
            O => \N__2576\,
            I => \myClockArea_timeout_counter_value_7\
        );

    \I__364\ : InMux
    port map (
            O => \N__2571\,
            I => \N__2567\
        );

    \I__363\ : InMux
    port map (
            O => \N__2570\,
            I => \N__2564\
        );

    \I__362\ : LocalMux
    port map (
            O => \N__2567\,
            I => \N__2561\
        );

    \I__361\ : LocalMux
    port map (
            O => \N__2564\,
            I => \myClockArea_timeout_counter_value_21\
        );

    \I__360\ : Odrv4
    port map (
            O => \N__2561\,
            I => \myClockArea_timeout_counter_value_21\
        );

    \I__359\ : CascadeMux
    port map (
            O => \N__2556\,
            I => \N__2552\
        );

    \I__358\ : InMux
    port map (
            O => \N__2555\,
            I => \N__2549\
        );

    \I__357\ : InMux
    port map (
            O => \N__2552\,
            I => \N__2546\
        );

    \I__356\ : LocalMux
    port map (
            O => \N__2549\,
            I => \ctrl_idcodeArea_shifter_5\
        );

    \I__355\ : LocalMux
    port map (
            O => \N__2546\,
            I => \ctrl_idcodeArea_shifter_5\
        );

    \I__354\ : CascadeMux
    port map (
            O => \N__2541\,
            I => \N__2537\
        );

    \I__353\ : InMux
    port map (
            O => \N__2540\,
            I => \N__2532\
        );

    \I__352\ : InMux
    port map (
            O => \N__2537\,
            I => \N__2532\
        );

    \I__351\ : LocalMux
    port map (
            O => \N__2532\,
            I => \ctrl_idcodeArea_shifter_7\
        );

    \I__350\ : CascadeMux
    port map (
            O => \N__2529\,
            I => \N__2525\
        );

    \I__349\ : InMux
    port map (
            O => \N__2528\,
            I => \N__2522\
        );

    \I__348\ : InMux
    port map (
            O => \N__2525\,
            I => \N__2519\
        );

    \I__347\ : LocalMux
    port map (
            O => \N__2522\,
            I => \ctrl_idcodeArea_shifter_6\
        );

    \I__346\ : LocalMux
    port map (
            O => \N__2519\,
            I => \ctrl_idcodeArea_shifter_6\
        );

    \I__345\ : InMux
    port map (
            O => \N__2514\,
            I => \N__2497\
        );

    \I__344\ : InMux
    port map (
            O => \N__2513\,
            I => \N__2497\
        );

    \I__343\ : InMux
    port map (
            O => \N__2512\,
            I => \N__2497\
        );

    \I__342\ : InMux
    port map (
            O => \N__2511\,
            I => \N__2497\
        );

    \I__341\ : InMux
    port map (
            O => \N__2510\,
            I => \N__2497\
        );

    \I__340\ : InMux
    port map (
            O => \N__2509\,
            I => \N__2492\
        );

    \I__339\ : InMux
    port map (
            O => \N__2508\,
            I => \N__2492\
        );

    \I__338\ : LocalMux
    port map (
            O => \N__2497\,
            I => n2045
        );

    \I__337\ : LocalMux
    port map (
            O => \N__2492\,
            I => n2045
        );

    \I__336\ : CascadeMux
    port map (
            O => \N__2487\,
            I => \N__2483\
        );

    \I__335\ : InMux
    port map (
            O => \N__2486\,
            I => \N__2480\
        );

    \I__334\ : InMux
    port map (
            O => \N__2483\,
            I => \N__2477\
        );

    \I__333\ : LocalMux
    port map (
            O => \N__2480\,
            I => \ctrl_idcodeArea_shifter_8\
        );

    \I__332\ : LocalMux
    port map (
            O => \N__2477\,
            I => \ctrl_idcodeArea_shifter_8\
        );

    \I__331\ : InMux
    port map (
            O => \N__2472\,
            I => \N__2469\
        );

    \I__330\ : LocalMux
    port map (
            O => \N__2469\,
            I => n2140
        );

    \I__329\ : CascadeMux
    port map (
            O => \N__2466\,
            I => \n9_cascade_\
        );

    \I__328\ : InMux
    port map (
            O => \N__2463\,
            I => \N__2460\
        );

    \I__327\ : LocalMux
    port map (
            O => \N__2460\,
            I => n2191
        );

    \I__326\ : InMux
    port map (
            O => \N__2457\,
            I => \N__2453\
        );

    \I__325\ : InMux
    port map (
            O => \N__2456\,
            I => \N__2450\
        );

    \I__324\ : LocalMux
    port map (
            O => \N__2453\,
            I => \ctrl_idcodeArea_shifter_25\
        );

    \I__323\ : LocalMux
    port map (
            O => \N__2450\,
            I => \ctrl_idcodeArea_shifter_25\
        );

    \I__322\ : InMux
    port map (
            O => \N__2445\,
            I => \N__2442\
        );

    \I__321\ : LocalMux
    port map (
            O => \N__2442\,
            I => n6
        );

    \I__320\ : InMux
    port map (
            O => \N__2439\,
            I => \N__2435\
        );

    \I__319\ : InMux
    port map (
            O => \N__2438\,
            I => \N__2432\
        );

    \I__318\ : LocalMux
    port map (
            O => \N__2435\,
            I => n1293
        );

    \I__317\ : LocalMux
    port map (
            O => \N__2432\,
            I => n1293
        );

    \I__316\ : CascadeMux
    port map (
            O => \N__2427\,
            I => \n1582_cascade_\
        );

    \I__315\ : InMux
    port map (
            O => \N__2424\,
            I => \N__2420\
        );

    \I__314\ : InMux
    port map (
            O => \N__2423\,
            I => \N__2417\
        );

    \I__313\ : LocalMux
    port map (
            O => \N__2420\,
            I => n2119
        );

    \I__312\ : LocalMux
    port map (
            O => \N__2417\,
            I => n2119
        );

    \I__311\ : InMux
    port map (
            O => \N__2412\,
            I => \N__2406\
        );

    \I__310\ : InMux
    port map (
            O => \N__2411\,
            I => \N__2406\
        );

    \I__309\ : LocalMux
    port map (
            O => \N__2406\,
            I => \ctrl_idcodeArea_shifter_24\
        );

    \I__308\ : CascadeMux
    port map (
            O => \N__2403\,
            I => \n2178_cascade_\
        );

    \I__307\ : InMux
    port map (
            O => \N__2400\,
            I => \N__2394\
        );

    \I__306\ : InMux
    port map (
            O => \N__2399\,
            I => \N__2394\
        );

    \I__305\ : LocalMux
    port map (
            O => \N__2394\,
            I => \ctrl_idcodeArea_shifter_23\
        );

    \I__304\ : CascadeMux
    port map (
            O => \N__2391\,
            I => \n1313_cascade_\
        );

    \I__303\ : InMux
    port map (
            O => \N__2388\,
            I => \N__2385\
        );

    \I__302\ : LocalMux
    port map (
            O => \N__2385\,
            I => \ctrl_tap_tdoUnbufferd_N_224\
        );

    \I__301\ : CascadeMux
    port map (
            O => \N__2382\,
            I => \N__2378\
        );

    \I__300\ : CascadeMux
    port map (
            O => \N__2381\,
            I => \N__2375\
        );

    \I__299\ : InMux
    port map (
            O => \N__2378\,
            I => \N__2372\
        );

    \I__298\ : InMux
    port map (
            O => \N__2375\,
            I => \N__2369\
        );

    \I__297\ : LocalMux
    port map (
            O => \N__2372\,
            I => \ctrl_idcodeArea_shifter_1\
        );

    \I__296\ : LocalMux
    port map (
            O => \N__2369\,
            I => \ctrl_idcodeArea_shifter_1\
        );

    \I__295\ : InMux
    port map (
            O => \N__2364\,
            I => \N__2360\
        );

    \I__294\ : InMux
    port map (
            O => \N__2363\,
            I => \N__2357\
        );

    \I__293\ : LocalMux
    port map (
            O => \N__2360\,
            I => \N__2354\
        );

    \I__292\ : LocalMux
    port map (
            O => \N__2357\,
            I => \ctrl_idcodeArea_shifter_0\
        );

    \I__291\ : Odrv4
    port map (
            O => \N__2354\,
            I => \ctrl_idcodeArea_shifter_0\
        );

    \I__290\ : CascadeMux
    port map (
            O => \N__2349\,
            I => \N__2345\
        );

    \I__289\ : InMux
    port map (
            O => \N__2348\,
            I => \N__2342\
        );

    \I__288\ : InMux
    port map (
            O => \N__2345\,
            I => \N__2339\
        );

    \I__287\ : LocalMux
    port map (
            O => \N__2342\,
            I => \ctrl_idcodeArea_shifter_29\
        );

    \I__286\ : LocalMux
    port map (
            O => \N__2339\,
            I => \ctrl_idcodeArea_shifter_29\
        );

    \I__285\ : CascadeMux
    port map (
            O => \N__2334\,
            I => \N__2331\
        );

    \I__284\ : InMux
    port map (
            O => \N__2331\,
            I => \N__2325\
        );

    \I__283\ : InMux
    port map (
            O => \N__2330\,
            I => \N__2325\
        );

    \I__282\ : LocalMux
    port map (
            O => \N__2325\,
            I => \ctrl_idcodeArea_shifter_28\
        );

    \I__281\ : CascadeMux
    port map (
            O => \N__2322\,
            I => \N__2319\
        );

    \I__280\ : InMux
    port map (
            O => \N__2319\,
            I => \N__2313\
        );

    \I__279\ : InMux
    port map (
            O => \N__2318\,
            I => \N__2313\
        );

    \I__278\ : LocalMux
    port map (
            O => \N__2313\,
            I => \ctrl_idcodeArea_shifter_27\
        );

    \I__277\ : CascadeMux
    port map (
            O => \N__2310\,
            I => \N__2307\
        );

    \I__276\ : InMux
    port map (
            O => \N__2307\,
            I => \N__2301\
        );

    \I__275\ : InMux
    port map (
            O => \N__2306\,
            I => \N__2301\
        );

    \I__274\ : LocalMux
    port map (
            O => \N__2301\,
            I => \ctrl_idcodeArea_shifter_26\
        );

    \I__273\ : InMux
    port map (
            O => \N__2298\,
            I => n2030
        );

    \I__272\ : InMux
    port map (
            O => \N__2295\,
            I => \N__2292\
        );

    \I__271\ : LocalMux
    port map (
            O => \N__2292\,
            I => n2116
        );

    \I__270\ : CascadeMux
    port map (
            O => \N__2289\,
            I => \n4_cascade_\
        );

    \I__269\ : CascadeMux
    port map (
            O => \N__2286\,
            I => \ctrl_tap_tdoUnbufferd_N_223_cascade_\
        );

    \I__268\ : IoInMux
    port map (
            O => \N__2283\,
            I => \N__2280\
        );

    \I__267\ : LocalMux
    port map (
            O => \N__2280\,
            I => \N__2277\
        );

    \I__266\ : IoSpan4Mux
    port map (
            O => \N__2277\,
            I => \N__2274\
        );

    \I__265\ : Odrv4
    port map (
            O => \N__2274\,
            I => \ctrl_tap_tdoUnbufferd\
        );

    \I__264\ : InMux
    port map (
            O => \N__2271\,
            I => \N__2261\
        );

    \I__263\ : InMux
    port map (
            O => \N__2270\,
            I => \N__2256\
        );

    \I__262\ : InMux
    port map (
            O => \N__2269\,
            I => \N__2256\
        );

    \I__261\ : InMux
    port map (
            O => \N__2268\,
            I => \N__2245\
        );

    \I__260\ : InMux
    port map (
            O => \N__2267\,
            I => \N__2245\
        );

    \I__259\ : InMux
    port map (
            O => \N__2266\,
            I => \N__2245\
        );

    \I__258\ : InMux
    port map (
            O => \N__2265\,
            I => \N__2245\
        );

    \I__257\ : InMux
    port map (
            O => \N__2264\,
            I => \N__2245\
        );

    \I__256\ : LocalMux
    port map (
            O => \N__2261\,
            I => n2146
        );

    \I__255\ : LocalMux
    port map (
            O => \N__2256\,
            I => n2146
        );

    \I__254\ : LocalMux
    port map (
            O => \N__2245\,
            I => n2146
        );

    \I__253\ : InMux
    port map (
            O => \N__2238\,
            I => n2021
        );

    \I__252\ : InMux
    port map (
            O => \N__2235\,
            I => n2022
        );

    \I__251\ : InMux
    port map (
            O => \N__2232\,
            I => n2023
        );

    \I__250\ : InMux
    port map (
            O => \N__2229\,
            I => \bfn_1_8_0_\
        );

    \I__249\ : InMux
    port map (
            O => \N__2226\,
            I => n2025
        );

    \I__248\ : InMux
    port map (
            O => \N__2223\,
            I => n2026
        );

    \I__247\ : InMux
    port map (
            O => \N__2220\,
            I => n2027
        );

    \I__246\ : InMux
    port map (
            O => \N__2217\,
            I => n2028
        );

    \I__245\ : InMux
    port map (
            O => \N__2214\,
            I => n2029
        );

    \I__244\ : InMux
    port map (
            O => \N__2211\,
            I => n2012
        );

    \I__243\ : InMux
    port map (
            O => \N__2208\,
            I => n2013
        );

    \I__242\ : InMux
    port map (
            O => \N__2205\,
            I => n2014
        );

    \I__241\ : InMux
    port map (
            O => \N__2202\,
            I => n2015
        );

    \I__240\ : InMux
    port map (
            O => \N__2199\,
            I => \bfn_1_7_0_\
        );

    \I__239\ : InMux
    port map (
            O => \N__2196\,
            I => n2017
        );

    \I__238\ : InMux
    port map (
            O => \N__2193\,
            I => n2018
        );

    \I__237\ : InMux
    port map (
            O => \N__2190\,
            I => n2019
        );

    \I__236\ : InMux
    port map (
            O => \N__2187\,
            I => n2020
        );

    \I__235\ : InMux
    port map (
            O => \N__2184\,
            I => \N__2181\
        );

    \I__234\ : LocalMux
    port map (
            O => \N__2181\,
            I => n1023
        );

    \I__233\ : InMux
    port map (
            O => \N__2178\,
            I => \N__2174\
        );

    \I__232\ : InMux
    port map (
            O => \N__2177\,
            I => \N__2171\
        );

    \I__231\ : LocalMux
    port map (
            O => \N__2174\,
            I => n1027
        );

    \I__230\ : LocalMux
    port map (
            O => \N__2171\,
            I => n1027
        );

    \I__229\ : InMux
    port map (
            O => \N__2166\,
            I => \N__2163\
        );

    \I__228\ : LocalMux
    port map (
            O => \N__2163\,
            I => n965
        );

    \I__227\ : InMux
    port map (
            O => \N__2160\,
            I => \N__2157\
        );

    \I__226\ : LocalMux
    port map (
            O => \N__2157\,
            I => n5
        );

    \I__225\ : CascadeMux
    port map (
            O => \N__2154\,
            I => \n5_cascade_\
        );

    \I__224\ : InMux
    port map (
            O => \N__2151\,
            I => \N__2148\
        );

    \I__223\ : LocalMux
    port map (
            O => \N__2148\,
            I => n2201
        );

    \I__222\ : InMux
    port map (
            O => \N__2145\,
            I => \bfn_1_6_0_\
        );

    \I__221\ : InMux
    port map (
            O => \N__2142\,
            I => n2009
        );

    \I__220\ : InMux
    port map (
            O => \N__2139\,
            I => n2010
        );

    \I__219\ : InMux
    port map (
            O => \N__2136\,
            I => n2011
        );

    \I__218\ : CascadeMux
    port map (
            O => \N__2133\,
            I => \n2188_cascade_\
        );

    \I__217\ : CascadeMux
    port map (
            O => \N__2130\,
            I => \n2235_cascade_\
        );

    \I__216\ : CascadeMux
    port map (
            O => \N__2127\,
            I => \n2202_cascade_\
        );

    \I__215\ : CascadeMux
    port map (
            O => \N__2124\,
            I => \N__2121\
        );

    \I__214\ : InMux
    port map (
            O => \N__2121\,
            I => \N__2118\
        );

    \I__213\ : LocalMux
    port map (
            O => \N__2118\,
            I => \N__2115\
        );

    \I__212\ : Odrv12
    port map (
            O => \N__2115\,
            I => n2211
        );

    \I__211\ : InMux
    port map (
            O => \N__2112\,
            I => \N__2109\
        );

    \I__210\ : LocalMux
    port map (
            O => \N__2109\,
            I => n962
        );

    \I__209\ : InMux
    port map (
            O => \N__2106\,
            I => \N__2103\
        );

    \I__208\ : LocalMux
    port map (
            O => \N__2103\,
            I => n1025
        );

    \I__207\ : CascadeMux
    port map (
            O => \N__2100\,
            I => \n1025_cascade_\
        );

    \I__206\ : CascadeMux
    port map (
            O => \N__2097\,
            I => \n960_cascade_\
        );

    \I__205\ : InMux
    port map (
            O => \N__2094\,
            I => \N__2091\
        );

    \I__204\ : LocalMux
    port map (
            O => \N__2091\,
            I => n2194
        );

    \I__203\ : CascadeMux
    port map (
            O => \N__2088\,
            I => \N__2085\
        );

    \I__202\ : InMux
    port map (
            O => \N__2085\,
            I => \N__2082\
        );

    \I__201\ : LocalMux
    port map (
            O => \N__2082\,
            I => n1828
        );

    \I__200\ : CascadeMux
    port map (
            O => \N__2079\,
            I => \n2045_cascade_\
        );

    \I__199\ : CascadeMux
    port map (
            O => \N__2076\,
            I => \N__2072\
        );

    \I__198\ : InMux
    port map (
            O => \N__2075\,
            I => \N__2067\
        );

    \I__197\ : InMux
    port map (
            O => \N__2072\,
            I => \N__2067\
        );

    \I__196\ : LocalMux
    port map (
            O => \N__2067\,
            I => \ctrl_idcodeArea_shifter_4\
        );

    \I__195\ : CascadeMux
    port map (
            O => \N__2064\,
            I => \N__2060\
        );

    \I__194\ : InMux
    port map (
            O => \N__2063\,
            I => \N__2057\
        );

    \I__193\ : InMux
    port map (
            O => \N__2060\,
            I => \N__2054\
        );

    \I__192\ : LocalMux
    port map (
            O => \N__2057\,
            I => \ctrl_idcodeArea_shifter_3\
        );

    \I__191\ : LocalMux
    port map (
            O => \N__2054\,
            I => \ctrl_idcodeArea_shifter_3\
        );

    \I__190\ : InMux
    port map (
            O => \N__2049\,
            I => \N__2043\
        );

    \I__189\ : InMux
    port map (
            O => \N__2048\,
            I => \N__2043\
        );

    \I__188\ : LocalMux
    port map (
            O => \N__2043\,
            I => \ctrl_idcodeArea_shifter_30\
        );

    \I__187\ : CascadeMux
    port map (
            O => \N__2040\,
            I => \n1854_cascade_\
        );

    \I__186\ : CascadeMux
    port map (
            O => \N__2037\,
            I => \n9_adj_2_cascade_\
        );

    \I__185\ : InMux
    port map (
            O => \N__2034\,
            I => \N__2031\
        );

    \I__184\ : LocalMux
    port map (
            O => \N__2031\,
            I => n8
        );

    \I__183\ : InMux
    port map (
            O => \N__2028\,
            I => \N__2025\
        );

    \I__182\ : LocalMux
    port map (
            O => \N__2025\,
            I => n12
        );

    \I__181\ : CascadeMux
    port map (
            O => \N__2022\,
            I => \n2_cascade_\
        );

    \I__180\ : InMux
    port map (
            O => \N__2019\,
            I => \N__2013\
        );

    \I__179\ : InMux
    port map (
            O => \N__2018\,
            I => \N__2013\
        );

    \I__178\ : LocalMux
    port map (
            O => \N__2013\,
            I => \ctrl_idcodeArea_shifter_2\
        );

    \I__177\ : CascadeMux
    port map (
            O => \N__2010\,
            I => \n12_cascade_\
        );

    \I__176\ : InMux
    port map (
            O => \N__2007\,
            I => \N__2004\
        );

    \I__175\ : LocalMux
    port map (
            O => \N__2004\,
            I => n1307
        );

    \I__174\ : CascadeMux
    port map (
            O => \N__2001\,
            I => \n2116_cascade_\
        );

    \I__173\ : IoInMux
    port map (
            O => \N__1998\,
            I => \N__1995\
        );

    \I__172\ : LocalMux
    port map (
            O => \N__1995\,
            I => \N__1992\
        );

    \I__171\ : Span4Mux_s3_h
    port map (
            O => \N__1992\,
            I => \N__1989\
        );

    \I__170\ : Sp12to4
    port map (
            O => \N__1989\,
            I => \N__1986\
        );

    \I__169\ : Odrv12
    port map (
            O => \N__1986\,
            I => io_jtag_tck_pad_gb_input
        );

    \IN_MUX_bfv_1_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_6_0_\
        );

    \IN_MUX_bfv_1_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n2016,
            carryinitout => \bfn_1_7_0_\
        );

    \IN_MUX_bfv_1_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n2024,
            carryinitout => \bfn_1_8_0_\
        );

    \io_jtag_tck_pad_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__1998\,
            GLOBALBUFFEROUTPUT => io_jtag_tck_c
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \i1_2_lut_adj_4_LC_1_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011101110"
        )
    port map (
            in0 => \N__3291\,
            in1 => \N__3186\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => n1307,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_tap_instruction_i1_LC_1_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100000000000"
        )
    port map (
            in0 => \N__3430\,
            in1 => \N__2269\,
            in2 => \N__3153\,
            in3 => \N__4921\,
            lcout => ctrl_tap_instruction_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4707\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \equal_312_i15_2_lut_LC_1_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3352\,
            in2 => \_gnd_net_\,
            in3 => \N__3334\,
            lcout => n12,
            ltout => \n12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_6_LC_1_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__3243\,
            in1 => \N__3396\,
            in2 => \N__2010\,
            in3 => \N__2007\,
            lcout => n2116,
            ltout => \n2116_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_adj_5_LC_1_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3429\,
            in2 => \N__2001\,
            in3 => \N__3126\,
            lcout => n15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_2_lut_3_lut_LC_1_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111010"
        )
    port map (
            in0 => \N__3187\,
            in1 => \_gnd_net_\,
            in2 => \N__3251\,
            in3 => \N__3292\,
            lcout => n8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_tap_instruction_i6_LC_1_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010100000100000"
        )
    port map (
            in0 => \N__4920\,
            in1 => \N__2271\,
            in2 => \N__3171\,
            in3 => \N__3188\,
            lcout => ctrl_tap_instruction_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4707\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_tap_instruction_i5_LC_1_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100000000000"
        )
    port map (
            in0 => \N__3335\,
            in1 => \N__2270\,
            in2 => \N__3321\,
            in3 => \N__4922\,
            lcout => ctrl_tap_instruction_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4707\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1047_2_lut_LC_1_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__3431\,
            in1 => \N__3127\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => n1828,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i20_3_lut_3_lut_LC_1_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010110101010"
        )
    port map (
            in0 => \N__3870\,
            in1 => \_gnd_net_\,
            in2 => \N__4214\,
            in3 => \N__3683\,
            lcout => OPEN,
            ltout => \n9_adj_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1424_3_lut_LC_1_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3937\,
            in2 => \N__2037\,
            in3 => \N__4076\,
            lcout => n2211,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_idcodeArea_shifter_i2_LC_1_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110000000000"
        )
    port map (
            in0 => \N__2018\,
            in1 => \N__2063\,
            in2 => \N__5082\,
            in3 => \N__4866\,
            lcout => \ctrl_idcodeArea_shifter_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4705\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_1_LC_1_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4184\,
            in2 => \_gnd_net_\,
            in3 => \N__3869\,
            lcout => OPEN,
            ltout => \n2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i5_4_lut_LC_1_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111111111"
        )
    port map (
            in0 => \N__2034\,
            in1 => \N__2028\,
            in2 => \N__2022\,
            in3 => \N__3397\,
            lcout => n1293,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1343_2_lut_3_lut_LC_1_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__3684\,
            in1 => \N__4188\,
            in2 => \_gnd_net_\,
            in3 => \N__3871\,
            lcout => n2146,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_idcodeArea_shifter_i1_LC_1_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010001000"
        )
    port map (
            in0 => \N__2019\,
            in1 => \N__4865\,
            in2 => \N__2381\,
            in3 => \N__5078\,
            lcout => \ctrl_idcodeArea_shifter_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4705\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_idcodeArea_shifter_i4_LC_1_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010001000"
        )
    port map (
            in0 => \N__2555\,
            in1 => \N__4859\,
            in2 => \N__2076\,
            in3 => \N__5048\,
            lcout => \ctrl_idcodeArea_shifter_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4703\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i3_4_lut_LC_1_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111111111111"
        )
    port map (
            in0 => \N__2438\,
            in1 => \N__3659\,
            in2 => \N__2088\,
            in3 => \N__4052\,
            lcout => n2045,
            ltout => \n2045_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_ledsArea_store_i0_i7_LC_1_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__4392\,
            in1 => \_gnd_net_\,
            in2 => \N__2079\,
            in3 => \N__4408\,
            lcout => io_leds_c_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4703\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_idcodeArea_shifter_i3_LC_1_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010000000000"
        )
    port map (
            in0 => \N__5075\,
            in1 => \N__2075\,
            in2 => \N__2064\,
            in3 => \N__4915\,
            lcout => \ctrl_idcodeArea_shifter_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4703\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_idcodeArea_shifter_i29_LC_1_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010001000"
        )
    port map (
            in0 => \N__2049\,
            in1 => \N__4858\,
            in2 => \N__2349\,
            in3 => \N__5047\,
            lcout => \ctrl_idcodeArea_shifter_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4703\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_idcodeArea_shifter_i30_LC_1_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101000010000000"
        )
    port map (
            in0 => \N__5074\,
            in1 => \N__2048\,
            in2 => \N__4916\,
            in3 => \N__3717\,
            lcout => \ctrl_idcodeArea_shifter_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4703\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_210_i4_4_lut_4_lut_LC_1_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101001001010"
        )
    port map (
            in0 => \N__4053\,
            in1 => \N__4178\,
            in2 => \N__3973\,
            in3 => \N__3864\,
            lcout => n962,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_tap_fsm_state_3__I_0_i6_2_lut_LC_1_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3658\,
            in2 => \_gnd_net_\,
            in3 => \N__4051\,
            lcout => n6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1073_2_lut_LC_1_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__3962\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2106\,
            lcout => OPEN,
            ltout => \n1854_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1385_4_lut_LC_1_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101011001100"
        )
    port map (
            in0 => \N__2178\,
            in1 => \N__3780\,
            in2 => \N__2040\,
            in3 => \N__2751\,
            lcout => OPEN,
            ltout => \n2188_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_tap_fsm_state_i2_LC_1_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__2753\,
            in1 => \N__2723\,
            in2 => \N__2133\,
            in3 => \N__2151\,
            lcout => ctrl_tap_fsm_state_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4701\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1431_2_lut_LC_1_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__4182\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2750\,
            lcout => OPEN,
            ltout => \n2235_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_tap_fsm_state_i0_LC_1_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111101001100"
        )
    port map (
            in0 => \N__3961\,
            in1 => \N__2721\,
            in2 => \N__2130\,
            in3 => \N__2094\,
            lcout => ctrl_tap_fsm_state_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4701\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1427_2_lut_4_lut_LC_1_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111011001100"
        )
    port map (
            in0 => \N__2160\,
            in1 => \N__3963\,
            in2 => \N__4213\,
            in3 => \N__3863\,
            lcout => OPEN,
            ltout => \n2202_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_tap_fsm_state_i1_LC_1_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__2752\,
            in1 => \N__2722\,
            in2 => \N__2127\,
            in3 => \N__2463\,
            lcout => ctrl_tap_fsm_state_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4701\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_tap_fsm_state_i3_LC_1_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101100010"
        )
    port map (
            in0 => \N__2724\,
            in1 => \N__2754\,
            in2 => \N__2124\,
            in3 => \N__2112\,
            lcout => ctrl_tap_fsm_state_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4701\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_3_lut_4_lut_LC_1_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__4171\,
            in1 => \N__4063\,
            in2 => \N__3691\,
            in3 => \N__3854\,
            lcout => n1025,
            ltout => \n1025_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_209_i1_4_lut_LC_1_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101001110111"
        )
    port map (
            in0 => \N__3968\,
            in1 => \N__2184\,
            in2 => \N__2100\,
            in3 => \N__2177\,
            lcout => OPEN,
            ltout => \n960_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1391_3_lut_LC_1_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2166\,
            in2 => \N__2097\,
            in3 => \N__2748\,
            lcout => n2194,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i3_2_lut_3_lut_4_lut_LC_1_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__3855\,
            in1 => \N__4168\,
            in2 => \N__4083\,
            in3 => \N__3663\,
            lcout => n1023,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_4_lut_adj_2_LC_1_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000110000"
        )
    port map (
            in0 => \N__4169\,
            in1 => \N__4062\,
            in2 => \N__3690\,
            in3 => \N__3853\,
            lcout => n1027,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_210_i1_4_lut_LC_1_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000110000"
        )
    port map (
            in0 => \N__3856\,
            in1 => \N__4170\,
            in2 => \N__3975\,
            in3 => \N__4068\,
            lcout => n965,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_LC_1_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__3670\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4064\,
            lcout => n5,
            ltout => \n5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1411_2_lut_4_lut_LC_1_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011111"
        )
    port map (
            in0 => \N__3857\,
            in1 => \N__3972\,
            in2 => \N__2154\,
            in3 => \N__4172\,
            lcout => n2201,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \myClockArea_timeout_counter_value_313__i0_LC_1_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__2907\,
            in1 => \N__2664\,
            in2 => \_gnd_net_\,
            in3 => \N__2145\,
            lcout => \myClockArea_timeout_counter_value_0\,
            ltout => OPEN,
            carryin => \bfn_1_6_0_\,
            carryout => n2009,
            clk => \N__5216\,
            ce => 'H',
            sr => \N__3486\
        );

    \myClockArea_timeout_counter_value_313__i1_LC_1_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__2877\,
            in1 => \N__2691\,
            in2 => \_gnd_net_\,
            in3 => \N__2142\,
            lcout => \myClockArea_timeout_counter_value_1\,
            ltout => OPEN,
            carryin => n2009,
            carryout => n2010,
            clk => \N__5216\,
            ce => 'H',
            sr => \N__3486\
        );

    \myClockArea_timeout_counter_value_313__i2_LC_1_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__2908\,
            in1 => \N__2967\,
            in2 => \_gnd_net_\,
            in3 => \N__2139\,
            lcout => \myClockArea_timeout_counter_value_2\,
            ltout => OPEN,
            carryin => n2010,
            carryout => n2011,
            clk => \N__5216\,
            ce => 'H',
            sr => \N__3486\
        );

    \myClockArea_timeout_counter_value_313__i3_LC_1_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__2878\,
            in1 => \N__2703\,
            in2 => \_gnd_net_\,
            in3 => \N__2136\,
            lcout => \myClockArea_timeout_counter_value_3\,
            ltout => OPEN,
            carryin => n2011,
            carryout => n2012,
            clk => \N__5216\,
            ce => 'H',
            sr => \N__3486\
        );

    \myClockArea_timeout_counter_value_313__i4_LC_1_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__2909\,
            in1 => \N__3057\,
            in2 => \_gnd_net_\,
            in3 => \N__2211\,
            lcout => \myClockArea_timeout_counter_value_4\,
            ltout => OPEN,
            carryin => n2012,
            carryout => n2013,
            clk => \N__5216\,
            ce => 'H',
            sr => \N__3486\
        );

    \myClockArea_timeout_counter_value_313__i5_LC_1_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__2879\,
            in1 => \N__2678\,
            in2 => \_gnd_net_\,
            in3 => \N__2208\,
            lcout => \myClockArea_timeout_counter_value_5\,
            ltout => OPEN,
            carryin => n2013,
            carryout => n2014,
            clk => \N__5216\,
            ce => 'H',
            sr => \N__3486\
        );

    \myClockArea_timeout_counter_value_313__i6_LC_1_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__2910\,
            in1 => \N__3045\,
            in2 => \_gnd_net_\,
            in3 => \N__2205\,
            lcout => \myClockArea_timeout_counter_value_6\,
            ltout => OPEN,
            carryin => n2014,
            carryout => n2015,
            clk => \N__5216\,
            ce => 'H',
            sr => \N__3486\
        );

    \myClockArea_timeout_counter_value_313__i7_LC_1_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__2880\,
            in1 => \N__2583\,
            in2 => \_gnd_net_\,
            in3 => \N__2202\,
            lcout => \myClockArea_timeout_counter_value_7\,
            ltout => OPEN,
            carryin => n2015,
            carryout => n2016,
            clk => \N__5216\,
            ce => 'H',
            sr => \N__3486\
        );

    \myClockArea_timeout_counter_value_313__i8_LC_1_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__2906\,
            in1 => \N__2994\,
            in2 => \_gnd_net_\,
            in3 => \N__2199\,
            lcout => \myClockArea_timeout_counter_value_8\,
            ltout => OPEN,
            carryin => \bfn_1_7_0_\,
            carryout => n2017,
            clk => \N__5215\,
            ce => 'H',
            sr => \N__3463\
        );

    \myClockArea_timeout_counter_value_313__i9_LC_1_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__2873\,
            in1 => \N__2652\,
            in2 => \_gnd_net_\,
            in3 => \N__2196\,
            lcout => \myClockArea_timeout_counter_value_9\,
            ltout => OPEN,
            carryin => n2017,
            carryout => n2018,
            clk => \N__5215\,
            ce => 'H',
            sr => \N__3463\
        );

    \myClockArea_timeout_counter_value_313__i10_LC_1_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__2903\,
            in1 => \N__2981\,
            in2 => \_gnd_net_\,
            in3 => \N__2193\,
            lcout => \myClockArea_timeout_counter_value_10\,
            ltout => OPEN,
            carryin => n2018,
            carryout => n2019,
            clk => \N__5215\,
            ce => 'H',
            sr => \N__3463\
        );

    \myClockArea_timeout_counter_value_313__i11_LC_1_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__2870\,
            in1 => \N__2778\,
            in2 => \_gnd_net_\,
            in3 => \N__2190\,
            lcout => \myClockArea_timeout_counter_value_11\,
            ltout => OPEN,
            carryin => n2019,
            carryout => n2020,
            clk => \N__5215\,
            ce => 'H',
            sr => \N__3463\
        );

    \myClockArea_timeout_counter_value_313__i12_LC_1_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__2904\,
            in1 => \N__2624\,
            in2 => \_gnd_net_\,
            in3 => \N__2187\,
            lcout => \myClockArea_timeout_counter_value_12\,
            ltout => OPEN,
            carryin => n2020,
            carryout => n2021,
            clk => \N__5215\,
            ce => 'H',
            sr => \N__3463\
        );

    \myClockArea_timeout_counter_value_313__i13_LC_1_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__2871\,
            in1 => \N__2940\,
            in2 => \_gnd_net_\,
            in3 => \N__2238\,
            lcout => \myClockArea_timeout_counter_value_13\,
            ltout => OPEN,
            carryin => n2021,
            carryout => n2022,
            clk => \N__5215\,
            ce => 'H',
            sr => \N__3463\
        );

    \myClockArea_timeout_counter_value_313__i14_LC_1_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__2905\,
            in1 => \N__2610\,
            in2 => \_gnd_net_\,
            in3 => \N__2235\,
            lcout => \myClockArea_timeout_counter_value_14\,
            ltout => OPEN,
            carryin => n2022,
            carryout => n2023,
            clk => \N__5215\,
            ce => 'H',
            sr => \N__3463\
        );

    \myClockArea_timeout_counter_value_313__i15_LC_1_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__2872\,
            in1 => \N__2805\,
            in2 => \_gnd_net_\,
            in3 => \N__2232\,
            lcout => \myClockArea_timeout_counter_value_15\,
            ltout => OPEN,
            carryin => n2023,
            carryout => n2024,
            clk => \N__5215\,
            ce => 'H',
            sr => \N__3463\
        );

    \myClockArea_timeout_counter_value_313__i16_LC_1_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__2899\,
            in1 => \N__3018\,
            in2 => \_gnd_net_\,
            in3 => \N__2229\,
            lcout => \myClockArea_timeout_counter_value_16\,
            ltout => OPEN,
            carryin => \bfn_1_8_0_\,
            carryout => n2025,
            clk => \N__5213\,
            ce => 'H',
            sr => \N__3478\
        );

    \myClockArea_timeout_counter_value_313__i17_LC_1_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__2874\,
            in1 => \N__3006\,
            in2 => \_gnd_net_\,
            in3 => \N__2226\,
            lcout => \myClockArea_timeout_counter_value_17\,
            ltout => OPEN,
            carryin => n2025,
            carryout => n2026,
            clk => \N__5213\,
            ce => 'H',
            sr => \N__3478\
        );

    \myClockArea_timeout_counter_value_313__i18_LC_1_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__2900\,
            in1 => \N__2639\,
            in2 => \_gnd_net_\,
            in3 => \N__2223\,
            lcout => \myClockArea_timeout_counter_value_18\,
            ltout => OPEN,
            carryin => n2026,
            carryout => n2027,
            clk => \N__5213\,
            ce => 'H',
            sr => \N__3478\
        );

    \myClockArea_timeout_counter_value_313__i19_LC_1_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__2875\,
            in1 => \N__2817\,
            in2 => \_gnd_net_\,
            in3 => \N__2220\,
            lcout => \myClockArea_timeout_counter_value_19\,
            ltout => OPEN,
            carryin => n2027,
            carryout => n2028,
            clk => \N__5213\,
            ce => 'H',
            sr => \N__3478\
        );

    \myClockArea_timeout_counter_value_313__i20_LC_1_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__2901\,
            in1 => \N__2792\,
            in2 => \_gnd_net_\,
            in3 => \N__2217\,
            lcout => \myClockArea_timeout_counter_value_20\,
            ltout => OPEN,
            carryin => n2028,
            carryout => n2029,
            clk => \N__5213\,
            ce => 'H',
            sr => \N__3478\
        );

    \myClockArea_timeout_counter_value_313__i21_LC_1_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__2876\,
            in1 => \N__2570\,
            in2 => \_gnd_net_\,
            in3 => \N__2214\,
            lcout => \myClockArea_timeout_counter_value_21\,
            ltout => OPEN,
            carryin => n2029,
            carryout => n2030,
            clk => \N__5213\,
            ce => 'H',
            sr => \N__3478\
        );

    \myClockArea_timeout_counter_value_313__i22_LC_1_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__2902\,
            in1 => \N__3032\,
            in2 => \_gnd_net_\,
            in3 => \N__2298\,
            lcout => \myClockArea_timeout_counter_value_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5213\,
            ce => 'H',
            sr => \N__3478\
        );

    \ctrl_tap_instruction_i4_LC_2_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100100001000000"
        )
    port map (
            in0 => \N__2265\,
            in1 => \N__4927\,
            in2 => \N__3273\,
            in3 => \N__3360\,
            lcout => ctrl_tap_instruction_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4710\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_tap_instruction_i0_LC_2_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100010100000"
        )
    port map (
            in0 => \N__4923\,
            in1 => \N__3128\,
            in2 => \N__3099\,
            in3 => \N__2268\,
            lcout => ctrl_tap_instruction_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4710\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_8_LC_2_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4341\,
            in2 => \_gnd_net_\,
            in3 => \N__2295\,
            lcout => OPEN,
            ltout => \n4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i395_4_lut_LC_2_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000000010"
        )
    port map (
            in0 => \N__2364\,
            in1 => \N__2423\,
            in2 => \N__2289\,
            in3 => \N__2388\,
            lcout => OPEN,
            ltout => \ctrl_tap_tdoUnbufferd_N_223_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i398_4_lut_LC_2_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__3509\,
            in1 => \N__3761\,
            in2 => \N__2286\,
            in3 => \N__4342\,
            lcout => \ctrl_tap_tdoUnbufferd\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_tap_instruction_i3_LC_2_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010100000100000"
        )
    port map (
            in0 => \N__4924\,
            in1 => \N__2266\,
            in2 => \N__3225\,
            in3 => \N__3247\,
            lcout => ctrl_tap_instruction_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4710\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_tap_instruction_i2_LC_2_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110110011"
        )
    port map (
            in0 => \N__2264\,
            in1 => \N__4926\,
            in2 => \N__3405\,
            in3 => \N__3375\,
            lcout => ctrl_tap_instruction_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4710\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_tap_instruction_i7_LC_2_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010001000"
        )
    port map (
            in0 => \N__4925\,
            in1 => \N__3207\,
            in2 => \N__3300\,
            in3 => \N__2267\,
            lcout => ctrl_tap_instruction_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4710\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_LC_2_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__4183\,
            in1 => \N__4072\,
            in2 => \_gnd_net_\,
            in3 => \N__3868\,
            lcout => OPEN,
            ltout => \n1313_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_tap_bypass_I_0_4_lut_LC_2_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110010101010"
        )
    port map (
            in0 => \N__5157\,
            in1 => \N__3092\,
            in2 => \N__2391\,
            in3 => \N__3682\,
            lcout => \ctrl_tap_tdoUnbufferd_N_224\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_idcodeArea_shifter_i25_LC_2_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011111111"
        )
    port map (
            in0 => \N__5039\,
            in1 => \N__2456\,
            in2 => \N__2310\,
            in3 => \N__4857\,
            lcout => \ctrl_idcodeArea_shifter_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4708\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_idcodeArea_shifter_i0_LC_2_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110101110101"
        )
    port map (
            in0 => \N__4854\,
            in1 => \N__5041\,
            in2 => \N__2382\,
            in3 => \N__2363\,
            lcout => \ctrl_idcodeArea_shifter_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4708\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_9_LC_2_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3125\,
            in2 => \_gnd_net_\,
            in3 => \N__3428\,
            lcout => n2119,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_idcodeArea_shifter_i28_LC_2_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010001000"
        )
    port map (
            in0 => \N__4856\,
            in1 => \N__2348\,
            in2 => \N__2334\,
            in3 => \N__5043\,
            lcout => \ctrl_idcodeArea_shifter_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4708\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_idcodeArea_shifter_i27_LC_2_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101000010000000"
        )
    port map (
            in0 => \N__5040\,
            in1 => \N__2318\,
            in2 => \N__4919\,
            in3 => \N__2330\,
            lcout => \ctrl_idcodeArea_shifter_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4708\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_idcodeArea_shifter_i26_LC_2_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110111110101"
        )
    port map (
            in0 => \N__4855\,
            in1 => \N__2306\,
            in2 => \N__2322\,
            in3 => \N__5042\,
            lcout => \ctrl_idcodeArea_shifter_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4708\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_idcodeArea_shifter_i22_LC_2_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111111001111"
        )
    port map (
            in0 => \N__3566\,
            in1 => \N__2400\,
            in2 => \N__4918\,
            in3 => \N__5038\,
            lcout => \ctrl_idcodeArea_shifter_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4706\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_tap_fsm_state_3__I_0_i7_2_lut_4_lut_LC_2_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__4146\,
            in1 => \N__4038\,
            in2 => \N__3681\,
            in3 => \N__3838\,
            lcout => n7_adj_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_ledsArea_store_i0_i5_LC_2_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__2509\,
            in1 => \N__4485\,
            in2 => \_gnd_net_\,
            in3 => \N__4496\,
            lcout => \ctrl_ledsArea_store_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4706\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_idcodeArea_shifter_i24_LC_2_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111101001111"
        )
    port map (
            in0 => \N__5037\,
            in1 => \N__2457\,
            in2 => \N__4917\,
            in3 => \N__2412\,
            lcout => \ctrl_idcodeArea_shifter_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4706\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_4_lut_adj_7_LC_2_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__3839\,
            in1 => \N__4147\,
            in2 => \N__4071\,
            in3 => \N__3649\,
            lcout => n1582,
            ltout => \n1582_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1375_4_lut_LC_2_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011100000"
        )
    port map (
            in0 => \N__2445\,
            in1 => \N__2439\,
            in2 => \N__2427\,
            in3 => \N__2424\,
            lcout => n2178,
            ltout => \n2178_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_idcodeArea_shifter_i23_LC_2_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101000000000"
        )
    port map (
            in0 => \N__2411\,
            in1 => \N__2399\,
            in2 => \N__2403\,
            in3 => \N__4870\,
            lcout => \ctrl_idcodeArea_shifter_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4706\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_ledsArea_store_i0_i1_LC_2_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__3532\,
            in1 => \N__2508\,
            in2 => \_gnd_net_\,
            in3 => \N__3510\,
            lcout => io_leds_c_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4706\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_idcodeArea_shifter_i7_LC_2_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010001000"
        )
    port map (
            in0 => \N__2486\,
            in1 => \N__4864\,
            in2 => \N__2541\,
            in3 => \N__5046\,
            lcout => \ctrl_idcodeArea_shifter_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4704\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_ledsArea_store_i0_i3_LC_2_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__2511\,
            in1 => \N__4575\,
            in2 => \_gnd_net_\,
            in3 => \N__4588\,
            lcout => io_leds_c_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4704\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_ledsArea_store_i0_i2_LC_2_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__4623\,
            in1 => \N__4636\,
            in2 => \_gnd_net_\,
            in3 => \N__2510\,
            lcout => io_leds_c_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4704\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_ledsArea_store_i0_i4_LC_2_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__2512\,
            in1 => \_gnd_net_\,
            in2 => \N__4524\,
            in3 => \N__4537\,
            lcout => io_leds_c_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4704\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_idcodeArea_shifter_i5_LC_2_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001110111011"
        )
    port map (
            in0 => \N__2528\,
            in1 => \N__4863\,
            in2 => \N__2556\,
            in3 => \N__5045\,
            lcout => \ctrl_idcodeArea_shifter_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4704\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_idcodeArea_shifter_i6_LC_2_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010000000000"
        )
    port map (
            in0 => \N__5044\,
            in1 => \N__2540\,
            in2 => \N__2529\,
            in3 => \N__4877\,
            lcout => \ctrl_idcodeArea_shifter_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4704\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_ledsArea_store_i0_i8_LC_2_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__4254\,
            in1 => \N__4306\,
            in2 => \_gnd_net_\,
            in3 => \N__2514\,
            lcout => io_leds_c_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4704\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_ledsArea_store_i0_i6_LC_2_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__2513\,
            in1 => \_gnd_net_\,
            in2 => \N__4434\,
            in3 => \N__4450\,
            lcout => io_leds_c_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4704\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1337_2_lut_LC_2_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3964\,
            in2 => \_gnd_net_\,
            in3 => \N__4065\,
            lcout => n2140,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_idcodeArea_shifter_i8_LC_2_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001110111011"
        )
    port map (
            in0 => \N__2597\,
            in1 => \N__4899\,
            in2 => \N__2487\,
            in3 => \N__5064\,
            lcout => \ctrl_idcodeArea_shifter_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4702\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i20_4_lut_3_lut_LC_2_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110001000"
        )
    port map (
            in0 => \N__4176\,
            in1 => \N__3677\,
            in2 => \_gnd_net_\,
            in3 => \N__3858\,
            lcout => OPEN,
            ltout => \n9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1388_4_lut_LC_2_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000000110011"
        )
    port map (
            in0 => \N__2472\,
            in1 => \N__2709\,
            in2 => \N__2466\,
            in3 => \N__2749\,
            lcout => n2191,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_LC_2_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001100110111"
        )
    port map (
            in0 => \N__4173\,
            in1 => \N__4066\,
            in2 => \N__3692\,
            in3 => \N__3859\,
            lcout => n12_adj_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i988_4_lut_4_lut_LC_2_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000000000001"
        )
    port map (
            in0 => \N__3861\,
            in1 => \N__4177\,
            in2 => \N__3694\,
            in3 => \N__4070\,
            lcout => n1769,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_4_lut_LC_2_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111111111"
        )
    port map (
            in0 => \N__4175\,
            in1 => \N__4067\,
            in2 => \N__3693\,
            in3 => \N__3862\,
            lcout => n7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_210_i2_4_lut_LC_2_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__3860\,
            in1 => \N__4174\,
            in2 => \N__3974\,
            in3 => \N__4069\,
            lcout => n1864,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1361_4_lut_LC_2_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__2702\,
            in1 => \N__2690\,
            in2 => \N__2679\,
            in3 => \N__2663\,
            lcout => n2164,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i5_4_lut_adj_3_LC_2_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__2651\,
            in1 => \N__2640\,
            in2 => \N__2625\,
            in3 => \N__2609\,
            lcout => n13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_idcodeArea_shifter_i9_LC_2_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010111011101"
        )
    port map (
            in0 => \N__4897\,
            in1 => \N__3066\,
            in2 => \N__2598\,
            in3 => \N__5063\,
            lcout => \ctrl_idcodeArea_shifter_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4700\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_idcodeArea_shifter_i11_LC_2_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100000000000"
        )
    port map (
            in0 => \N__5061\,
            in1 => \N__3074\,
            in2 => \N__5112\,
            in3 => \N__4898\,
            lcout => \ctrl_idcodeArea_shifter_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4700\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i3_2_lut_LC_2_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2582\,
            in2 => \_gnd_net_\,
            in3 => \N__2571\,
            lcout => n11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_idcodeArea_shifter_i10_LC_2_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100010100000"
        )
    port map (
            in0 => \N__4896\,
            in1 => \N__3065\,
            in2 => \N__3078\,
            in3 => \N__5062\,
            lcout => \ctrl_idcodeArea_shifter_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4700\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1373_4_lut_LC_2_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__3056\,
            in1 => \N__3044\,
            in2 => \N__3033\,
            in3 => \N__3017\,
            lcout => n2176,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1357_4_lut_LC_2_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__3005\,
            in1 => \N__2993\,
            in2 => \N__2982\,
            in3 => \N__2966\,
            lcout => OPEN,
            ltout => \n2160_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1379_4_lut_LC_2_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__2955\,
            in1 => \N__2766\,
            in2 => \N__2949\,
            in3 => \N__2946\,
            lcout => OPEN,
            ltout => \n2182_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i7_4_lut_LC_2_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__2939\,
            in1 => \N__2928\,
            in2 => \N__2922\,
            in3 => \N__2919\,
            lcout => n2113,
            ltout => \n2113_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i990_2_lut_LC_2_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2913\,
            in3 => \N__5261\,
            lcout => n1771,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1359_4_lut_LC_2_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__2816\,
            in1 => \N__2804\,
            in2 => \N__2793\,
            in3 => \N__2777\,
            lcout => n2162,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \myClockArea_timeout_state_88_LC_2_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5257\,
            in2 => \_gnd_net_\,
            in3 => \N__2760\,
            lcout => \myClockArea_timeout_state\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5214\,
            ce => 'H',
            sr => \N__3485\
        );

    \ctrl_tap_instructionShift_i0_i1_LC_4_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__4217\,
            in1 => \N__3371\,
            in2 => \_gnd_net_\,
            in3 => \N__3435\,
            lcout => \ctrl_tap_instructionShift_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4714\,
            ce => \N__3594\,
            sr => \_gnd_net_\
        );

    \ctrl_tap_instructionShift_i0_i2_LC_4_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__3218\,
            in1 => \N__3404\,
            in2 => \_gnd_net_\,
            in3 => \N__4222\,
            lcout => \ctrl_tap_instructionShift_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4714\,
            ce => \N__3594\,
            sr => \_gnd_net_\
        );

    \ctrl_tap_instructionShift_i0_i4_LC_4_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__4218\,
            in1 => \N__3311\,
            in2 => \_gnd_net_\,
            in3 => \N__3359\,
            lcout => \ctrl_tap_instructionShift_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4714\,
            ce => \N__3594\,
            sr => \_gnd_net_\
        );

    \ctrl_tap_instructionShift_i0_i5_LC_4_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__3164\,
            in1 => \N__4221\,
            in2 => \_gnd_net_\,
            in3 => \N__3339\,
            lcout => \ctrl_tap_instructionShift_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4714\,
            ce => \N__3594\,
            sr => \_gnd_net_\
        );

    \ctrl_tap_instructionShift_i0_i7_LC_4_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__4220\,
            in1 => \N__5181\,
            in2 => \_gnd_net_\,
            in3 => \N__3299\,
            lcout => \ctrl_tap_instructionShift_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4714\,
            ce => \N__3594\,
            sr => \_gnd_net_\
        );

    \ctrl_tap_instructionShift_i0_i3_LC_4_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__3263\,
            in1 => \N__3252\,
            in2 => \_gnd_net_\,
            in3 => \N__4223\,
            lcout => \ctrl_tap_instructionShift_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4714\,
            ce => \N__3594\,
            sr => \_gnd_net_\
        );

    \ctrl_tap_instructionShift_i0_i6_LC_4_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__4219\,
            in1 => \N__3203\,
            in2 => \_gnd_net_\,
            in3 => \N__3192\,
            lcout => \ctrl_tap_instructionShift_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4714\,
            ce => \N__3594\,
            sr => \_gnd_net_\
        );

    \ctrl_tap_instructionShift_i0_i0_LC_4_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__3146\,
            in1 => \N__3135\,
            in2 => \_gnd_net_\,
            in3 => \N__4224\,
            lcout => \ctrl_tap_instructionShift_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4712\,
            ce => \N__3590\,
            sr => \_gnd_net_\
        );

    \i1436_2_lut_3_lut_4_lut_LC_4_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__4086\,
            in1 => \N__3768\,
            in2 => \N__3702\,
            in3 => \N__3881\,
            lcout => n1353,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_idcodeArea_shifter_i18_LC_4_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101111110001111"
        )
    port map (
            in0 => \N__5049\,
            in1 => \N__3746\,
            in2 => \N__4928\,
            in3 => \N__3726\,
            lcout => \ctrl_idcodeArea_shifter_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4711\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_idcodeArea_shifter_i17_LC_4_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011000000"
        )
    port map (
            in0 => \N__5144\,
            in1 => \N__4900\,
            in2 => \N__3750\,
            in3 => \N__5053\,
            lcout => \ctrl_idcodeArea_shifter_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4711\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_idcodeArea_shifter_i20_LC_4_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010000000000"
        )
    port map (
            in0 => \N__5050\,
            in1 => \N__3555\,
            in2 => \N__3738\,
            in3 => \N__4911\,
            lcout => \ctrl_idcodeArea_shifter_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4711\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_idcodeArea_shifter_i19_LC_4_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110000000000"
        )
    port map (
            in0 => \N__3725\,
            in1 => \N__3737\,
            in2 => \N__5077\,
            in3 => \N__4904\,
            lcout => \ctrl_idcodeArea_shifter_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4711\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_idcodeArea_shifter_i31_LC_4_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011111111"
        )
    port map (
            in0 => \N__5052\,
            in1 => \N__3716\,
            in2 => \N__5195\,
            in3 => \N__4913\,
            lcout => \ctrl_idcodeArea_shifter_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4711\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_4_lut_LC_4_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000010000"
        )
    port map (
            in0 => \N__4216\,
            in1 => \N__4085\,
            in2 => \N__3701\,
            in3 => \N__3882\,
            lcout => n1067,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_idcodeArea_shifter_i21_LC_4_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011111111"
        )
    port map (
            in0 => \N__5051\,
            in1 => \N__3554\,
            in2 => \N__3573\,
            in3 => \N__4912\,
            lcout => \ctrl_idcodeArea_shifter_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4711\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_ledsArea_shifter_i0_i0_LC_4_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__3539\,
            in1 => \N__4283\,
            in2 => \N__4622\,
            in3 => \N__4365\,
            lcout => \ctrl_ledsArea_shifter_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4709\,
            ce => \N__4236\,
            sr => \_gnd_net_\
        );

    \ctrl_ledsArea_shifter_i0_i1_LC_4_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011100100"
        )
    port map (
            in0 => \N__4361\,
            in1 => \N__4571\,
            in2 => \N__4649\,
            in3 => \N__4287\,
            lcout => \ctrl_ledsArea_shifter_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4709\,
            ce => \N__4236\,
            sr => \_gnd_net_\
        );

    \ctrl_ledsArea_shifter_i0_i2_LC_4_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__4595\,
            in1 => \N__4284\,
            in2 => \N__4520\,
            in3 => \N__4366\,
            lcout => \ctrl_ledsArea_shifter_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4709\,
            ce => \N__4236\,
            sr => \_gnd_net_\
        );

    \ctrl_ledsArea_shifter_i0_i3_LC_4_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__4362\,
            in1 => \N__4544\,
            in2 => \N__4481\,
            in3 => \N__4288\,
            lcout => \ctrl_ledsArea_shifter_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4709\,
            ce => \N__4236\,
            sr => \_gnd_net_\
        );

    \ctrl_ledsArea_shifter_i0_i4_LC_4_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010111100100000"
        )
    port map (
            in0 => \N__4503\,
            in1 => \N__4285\,
            in2 => \N__4371\,
            in3 => \N__4427\,
            lcout => \ctrl_ledsArea_shifter_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4709\,
            ce => \N__4236\,
            sr => \_gnd_net_\
        );

    \ctrl_ledsArea_shifter_i0_i5_LC_4_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__4363\,
            in1 => \N__4457\,
            in2 => \N__4388\,
            in3 => \N__4289\,
            lcout => \ctrl_ledsArea_shifter_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4709\,
            ce => \N__4236\,
            sr => \_gnd_net_\
        );

    \ctrl_ledsArea_shifter_i0_i6_LC_4_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__4416\,
            in1 => \N__4286\,
            in2 => \N__4253\,
            in3 => \N__4367\,
            lcout => \ctrl_ledsArea_shifter_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4709\,
            ce => \N__4236\,
            sr => \_gnd_net_\
        );

    \ctrl_ledsArea_shifter_i0_i7_LC_4_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__4364\,
            in1 => \N__4313\,
            in2 => \N__5196\,
            in3 => \N__4290\,
            lcout => \ctrl_ledsArea_shifter_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4709\,
            ce => \N__4236\,
            sr => \_gnd_net_\
        );

    \mux_210_i3_4_lut_4_lut_LC_4_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101001100010011"
        )
    port map (
            in0 => \N__4215\,
            in1 => \N__4084\,
            in2 => \N__3933\,
            in3 => \N__3880\,
            lcout => n963,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \myClockArea_toggle_90_LC_4_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5228\,
            in2 => \_gnd_net_\,
            in3 => \N__5262\,
            lcout => io_leds_c_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5217\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_tap_bypass_81_LC_5_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5185\,
            lcout => ctrl_tap_bypass,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4715\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_idcodeArea_shifter_i14_LC_5_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011111111"
        )
    port map (
            in0 => \N__5055\,
            in1 => \N__5132\,
            in2 => \N__4728\,
            in3 => \N__4914\,
            lcout => \ctrl_idcodeArea_shifter_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4713\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_idcodeArea_shifter_i16_LC_5_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101111110011"
        )
    port map (
            in0 => \N__5090\,
            in1 => \N__4906\,
            in2 => \N__5148\,
            in3 => \N__5057\,
            lcout => \ctrl_idcodeArea_shifter_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4713\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_idcodeArea_shifter_i13_LC_5_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101000010000000"
        )
    port map (
            in0 => \N__5054\,
            in1 => \N__5120\,
            in2 => \N__4929\,
            in3 => \N__5133\,
            lcout => \ctrl_idcodeArea_shifter_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4713\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_idcodeArea_shifter_i12_LC_5_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011000000"
        )
    port map (
            in0 => \N__5102\,
            in1 => \N__4905\,
            in2 => \N__5124\,
            in3 => \N__5056\,
            lcout => \ctrl_idcodeArea_shifter_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4713\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_idcodeArea_shifter_i15_LC_5_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101000000000"
        )
    port map (
            in0 => \N__5091\,
            in1 => \N__4727\,
            in2 => \N__5076\,
            in3 => \N__4910\,
            lcout => \ctrl_idcodeArea_shifter_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4713\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
