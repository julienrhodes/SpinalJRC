// ******************************************************************************

// iCEcube Netlister

// Version:            2017.08.27940

// Build Date:         Sep 12 2017 08:25:46

// File Generated:     May 5 2020 16:11:55

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "MyTopLevel" view "INTERFACE"

module MyTopLevel (
    io_leds,
    io_jtag_tms,
    io_jtag_tdo,
    io_jtag_tdi,
    io_jtag_tck,
    global_reset,
    global_clk);

    output [7:0] io_leds;
    input io_jtag_tms;
    output io_jtag_tdo;
    input io_jtag_tdi;
    input io_jtag_tck;
    input global_reset;
    input global_clk;

    wire N__4910;
    wire N__4909;
    wire N__4908;
    wire N__4899;
    wire N__4898;
    wire N__4897;
    wire N__4890;
    wire N__4889;
    wire N__4888;
    wire N__4881;
    wire N__4880;
    wire N__4879;
    wire N__4872;
    wire N__4871;
    wire N__4870;
    wire N__4863;
    wire N__4862;
    wire N__4861;
    wire N__4854;
    wire N__4853;
    wire N__4852;
    wire N__4845;
    wire N__4844;
    wire N__4843;
    wire N__4836;
    wire N__4835;
    wire N__4834;
    wire N__4827;
    wire N__4826;
    wire N__4825;
    wire N__4818;
    wire N__4817;
    wire N__4816;
    wire N__4809;
    wire N__4808;
    wire N__4807;
    wire N__4800;
    wire N__4799;
    wire N__4798;
    wire N__4791;
    wire N__4790;
    wire N__4789;
    wire N__4772;
    wire N__4769;
    wire N__4766;
    wire N__4763;
    wire N__4762;
    wire N__4759;
    wire N__4756;
    wire N__4755;
    wire N__4752;
    wire N__4749;
    wire N__4746;
    wire N__4739;
    wire N__4738;
    wire N__4735;
    wire N__4732;
    wire N__4729;
    wire N__4724;
    wire N__4721;
    wire N__4720;
    wire N__4717;
    wire N__4714;
    wire N__4709;
    wire N__4708;
    wire N__4705;
    wire N__4702;
    wire N__4697;
    wire N__4696;
    wire N__4693;
    wire N__4690;
    wire N__4687;
    wire N__4684;
    wire N__4681;
    wire N__4678;
    wire N__4677;
    wire N__4672;
    wire N__4669;
    wire N__4664;
    wire N__4663;
    wire N__4660;
    wire N__4657;
    wire N__4654;
    wire N__4651;
    wire N__4648;
    wire N__4643;
    wire N__4642;
    wire N__4639;
    wire N__4636;
    wire N__4633;
    wire N__4628;
    wire N__4627;
    wire N__4626;
    wire N__4625;
    wire N__4624;
    wire N__4619;
    wire N__4612;
    wire N__4607;
    wire N__4604;
    wire N__4601;
    wire N__4600;
    wire N__4597;
    wire N__4594;
    wire N__4591;
    wire N__4588;
    wire N__4583;
    wire N__4582;
    wire N__4579;
    wire N__4576;
    wire N__4571;
    wire N__4570;
    wire N__4567;
    wire N__4564;
    wire N__4561;
    wire N__4558;
    wire N__4557;
    wire N__4556;
    wire N__4555;
    wire N__4554;
    wire N__4553;
    wire N__4552;
    wire N__4551;
    wire N__4548;
    wire N__4545;
    wire N__4534;
    wire N__4529;
    wire N__4520;
    wire N__4517;
    wire N__4514;
    wire N__4513;
    wire N__4510;
    wire N__4507;
    wire N__4502;
    wire N__4499;
    wire N__4498;
    wire N__4497;
    wire N__4494;
    wire N__4491;
    wire N__4488;
    wire N__4485;
    wire N__4482;
    wire N__4479;
    wire N__4472;
    wire N__4471;
    wire N__4468;
    wire N__4465;
    wire N__4462;
    wire N__4457;
    wire N__4454;
    wire N__4451;
    wire N__4450;
    wire N__4449;
    wire N__4446;
    wire N__4443;
    wire N__4440;
    wire N__4433;
    wire N__4430;
    wire N__4429;
    wire N__4426;
    wire N__4423;
    wire N__4418;
    wire N__4417;
    wire N__4416;
    wire N__4415;
    wire N__4414;
    wire N__4411;
    wire N__4408;
    wire N__4405;
    wire N__4402;
    wire N__4401;
    wire N__4400;
    wire N__4397;
    wire N__4394;
    wire N__4393;
    wire N__4388;
    wire N__4385;
    wire N__4380;
    wire N__4377;
    wire N__4374;
    wire N__4371;
    wire N__4364;
    wire N__4355;
    wire N__4352;
    wire N__4351;
    wire N__4348;
    wire N__4345;
    wire N__4342;
    wire N__4339;
    wire N__4338;
    wire N__4335;
    wire N__4332;
    wire N__4329;
    wire N__4322;
    wire N__4321;
    wire N__4320;
    wire N__4319;
    wire N__4318;
    wire N__4317;
    wire N__4316;
    wire N__4315;
    wire N__4314;
    wire N__4313;
    wire N__4312;
    wire N__4311;
    wire N__4310;
    wire N__4309;
    wire N__4308;
    wire N__4307;
    wire N__4306;
    wire N__4305;
    wire N__4304;
    wire N__4265;
    wire N__4262;
    wire N__4259;
    wire N__4258;
    wire N__4255;
    wire N__4252;
    wire N__4247;
    wire N__4244;
    wire N__4241;
    wire N__4238;
    wire N__4235;
    wire N__4232;
    wire N__4231;
    wire N__4228;
    wire N__4227;
    wire N__4226;
    wire N__4223;
    wire N__4220;
    wire N__4215;
    wire N__4208;
    wire N__4205;
    wire N__4204;
    wire N__4203;
    wire N__4202;
    wire N__4201;
    wire N__4200;
    wire N__4199;
    wire N__4198;
    wire N__4195;
    wire N__4192;
    wire N__4189;
    wire N__4184;
    wire N__4181;
    wire N__4178;
    wire N__4175;
    wire N__4160;
    wire N__4157;
    wire N__4156;
    wire N__4155;
    wire N__4154;
    wire N__4153;
    wire N__4152;
    wire N__4145;
    wire N__4144;
    wire N__4143;
    wire N__4142;
    wire N__4141;
    wire N__4140;
    wire N__4137;
    wire N__4134;
    wire N__4131;
    wire N__4128;
    wire N__4125;
    wire N__4124;
    wire N__4123;
    wire N__4122;
    wire N__4121;
    wire N__4120;
    wire N__4117;
    wire N__4116;
    wire N__4115;
    wire N__4114;
    wire N__4113;
    wire N__4112;
    wire N__4111;
    wire N__4110;
    wire N__4107;
    wire N__4100;
    wire N__4095;
    wire N__4092;
    wire N__4083;
    wire N__4076;
    wire N__4067;
    wire N__4060;
    wire N__4043;
    wire N__4042;
    wire N__4041;
    wire N__4040;
    wire N__4039;
    wire N__4038;
    wire N__4037;
    wire N__4036;
    wire N__4035;
    wire N__4034;
    wire N__4033;
    wire N__4032;
    wire N__4029;
    wire N__4028;
    wire N__4027;
    wire N__4024;
    wire N__4023;
    wire N__4022;
    wire N__4021;
    wire N__4018;
    wire N__4017;
    wire N__4010;
    wire N__4007;
    wire N__4004;
    wire N__4001;
    wire N__3996;
    wire N__3987;
    wire N__3980;
    wire N__3973;
    wire N__3956;
    wire N__3955;
    wire N__3954;
    wire N__3953;
    wire N__3952;
    wire N__3951;
    wire N__3950;
    wire N__3949;
    wire N__3946;
    wire N__3945;
    wire N__3944;
    wire N__3943;
    wire N__3940;
    wire N__3939;
    wire N__3934;
    wire N__3931;
    wire N__3926;
    wire N__3923;
    wire N__3920;
    wire N__3913;
    wire N__3912;
    wire N__3907;
    wire N__3900;
    wire N__3897;
    wire N__3892;
    wire N__3889;
    wire N__3886;
    wire N__3883;
    wire N__3880;
    wire N__3877;
    wire N__3874;
    wire N__3871;
    wire N__3868;
    wire N__3865;
    wire N__3860;
    wire N__3851;
    wire N__3850;
    wire N__3849;
    wire N__3848;
    wire N__3847;
    wire N__3844;
    wire N__3843;
    wire N__3842;
    wire N__3841;
    wire N__3840;
    wire N__3839;
    wire N__3838;
    wire N__3837;
    wire N__3836;
    wire N__3829;
    wire N__3826;
    wire N__3823;
    wire N__3822;
    wire N__3821;
    wire N__3820;
    wire N__3819;
    wire N__3818;
    wire N__3817;
    wire N__3816;
    wire N__3815;
    wire N__3814;
    wire N__3807;
    wire N__3804;
    wire N__3799;
    wire N__3794;
    wire N__3791;
    wire N__3786;
    wire N__3779;
    wire N__3774;
    wire N__3765;
    wire N__3746;
    wire N__3743;
    wire N__3740;
    wire N__3737;
    wire N__3734;
    wire N__3733;
    wire N__3732;
    wire N__3731;
    wire N__3730;
    wire N__3727;
    wire N__3726;
    wire N__3725;
    wire N__3724;
    wire N__3723;
    wire N__3722;
    wire N__3721;
    wire N__3720;
    wire N__3719;
    wire N__3716;
    wire N__3715;
    wire N__3712;
    wire N__3711;
    wire N__3708;
    wire N__3707;
    wire N__3706;
    wire N__3705;
    wire N__3704;
    wire N__3703;
    wire N__3700;
    wire N__3699;
    wire N__3698;
    wire N__3697;
    wire N__3694;
    wire N__3689;
    wire N__3680;
    wire N__3677;
    wire N__3672;
    wire N__3669;
    wire N__3664;
    wire N__3661;
    wire N__3656;
    wire N__3649;
    wire N__3644;
    wire N__3639;
    wire N__3614;
    wire N__3611;
    wire N__3608;
    wire N__3605;
    wire N__3602;
    wire N__3599;
    wire N__3596;
    wire N__3593;
    wire N__3590;
    wire N__3589;
    wire N__3586;
    wire N__3583;
    wire N__3580;
    wire N__3575;
    wire N__3572;
    wire N__3569;
    wire N__3566;
    wire N__3563;
    wire N__3560;
    wire N__3557;
    wire N__3554;
    wire N__3551;
    wire N__3550;
    wire N__3547;
    wire N__3544;
    wire N__3539;
    wire N__3538;
    wire N__3535;
    wire N__3532;
    wire N__3527;
    wire N__3524;
    wire N__3523;
    wire N__3522;
    wire N__3519;
    wire N__3516;
    wire N__3513;
    wire N__3512;
    wire N__3509;
    wire N__3506;
    wire N__3503;
    wire N__3500;
    wire N__3495;
    wire N__3490;
    wire N__3485;
    wire N__3484;
    wire N__3481;
    wire N__3478;
    wire N__3475;
    wire N__3470;
    wire N__3469;
    wire N__3466;
    wire N__3463;
    wire N__3460;
    wire N__3455;
    wire N__3454;
    wire N__3449;
    wire N__3446;
    wire N__3445;
    wire N__3442;
    wire N__3439;
    wire N__3436;
    wire N__3431;
    wire N__3430;
    wire N__3429;
    wire N__3428;
    wire N__3427;
    wire N__3426;
    wire N__3425;
    wire N__3424;
    wire N__3423;
    wire N__3422;
    wire N__3421;
    wire N__3420;
    wire N__3419;
    wire N__3418;
    wire N__3417;
    wire N__3416;
    wire N__3415;
    wire N__3414;
    wire N__3413;
    wire N__3412;
    wire N__3411;
    wire N__3410;
    wire N__3409;
    wire N__3408;
    wire N__3407;
    wire N__3406;
    wire N__3405;
    wire N__3404;
    wire N__3403;
    wire N__3402;
    wire N__3401;
    wire N__3400;
    wire N__3397;
    wire N__3388;
    wire N__3371;
    wire N__3360;
    wire N__3349;
    wire N__3332;
    wire N__3327;
    wire N__3314;
    wire N__3313;
    wire N__3310;
    wire N__3307;
    wire N__3302;
    wire N__3299;
    wire N__3298;
    wire N__3297;
    wire N__3296;
    wire N__3295;
    wire N__3294;
    wire N__3293;
    wire N__3292;
    wire N__3291;
    wire N__3290;
    wire N__3287;
    wire N__3286;
    wire N__3285;
    wire N__3282;
    wire N__3279;
    wire N__3278;
    wire N__3275;
    wire N__3272;
    wire N__3271;
    wire N__3270;
    wire N__3267;
    wire N__3266;
    wire N__3263;
    wire N__3260;
    wire N__3259;
    wire N__3250;
    wire N__3249;
    wire N__3248;
    wire N__3247;
    wire N__3246;
    wire N__3245;
    wire N__3244;
    wire N__3243;
    wire N__3242;
    wire N__3241;
    wire N__3240;
    wire N__3239;
    wire N__3238;
    wire N__3237;
    wire N__3220;
    wire N__3209;
    wire N__3208;
    wire N__3207;
    wire N__3206;
    wire N__3205;
    wire N__3204;
    wire N__3203;
    wire N__3200;
    wire N__3193;
    wire N__3188;
    wire N__3179;
    wire N__3170;
    wire N__3165;
    wire N__3160;
    wire N__3151;
    wire N__3134;
    wire N__3133;
    wire N__3130;
    wire N__3125;
    wire N__3122;
    wire N__3119;
    wire N__3118;
    wire N__3117;
    wire N__3116;
    wire N__3115;
    wire N__3114;
    wire N__3113;
    wire N__3112;
    wire N__3111;
    wire N__3110;
    wire N__3109;
    wire N__3108;
    wire N__3099;
    wire N__3098;
    wire N__3097;
    wire N__3096;
    wire N__3095;
    wire N__3094;
    wire N__3093;
    wire N__3092;
    wire N__3091;
    wire N__3090;
    wire N__3089;
    wire N__3088;
    wire N__3079;
    wire N__3070;
    wire N__3067;
    wire N__3058;
    wire N__3051;
    wire N__3042;
    wire N__3029;
    wire N__3028;
    wire N__3025;
    wire N__3022;
    wire N__3017;
    wire N__3016;
    wire N__3013;
    wire N__3010;
    wire N__3005;
    wire N__3002;
    wire N__2999;
    wire N__2998;
    wire N__2995;
    wire N__2992;
    wire N__2987;
    wire N__2986;
    wire N__2983;
    wire N__2980;
    wire N__2975;
    wire N__2974;
    wire N__2971;
    wire N__2968;
    wire N__2965;
    wire N__2960;
    wire N__2959;
    wire N__2956;
    wire N__2953;
    wire N__2948;
    wire N__2945;
    wire N__2942;
    wire N__2941;
    wire N__2938;
    wire N__2935;
    wire N__2930;
    wire N__2929;
    wire N__2926;
    wire N__2923;
    wire N__2918;
    wire N__2917;
    wire N__2914;
    wire N__2911;
    wire N__2908;
    wire N__2903;
    wire N__2902;
    wire N__2899;
    wire N__2896;
    wire N__2891;
    wire N__2888;
    wire N__2885;
    wire N__2884;
    wire N__2883;
    wire N__2880;
    wire N__2877;
    wire N__2874;
    wire N__2871;
    wire N__2864;
    wire N__2861;
    wire N__2860;
    wire N__2857;
    wire N__2854;
    wire N__2849;
    wire N__2848;
    wire N__2847;
    wire N__2846;
    wire N__2845;
    wire N__2834;
    wire N__2831;
    wire N__2828;
    wire N__2827;
    wire N__2822;
    wire N__2819;
    wire N__2818;
    wire N__2815;
    wire N__2810;
    wire N__2807;
    wire N__2804;
    wire N__2801;
    wire N__2800;
    wire N__2797;
    wire N__2796;
    wire N__2793;
    wire N__2790;
    wire N__2787;
    wire N__2784;
    wire N__2777;
    wire N__2776;
    wire N__2773;
    wire N__2770;
    wire N__2765;
    wire N__2764;
    wire N__2761;
    wire N__2758;
    wire N__2753;
    wire N__2752;
    wire N__2749;
    wire N__2746;
    wire N__2743;
    wire N__2738;
    wire N__2737;
    wire N__2734;
    wire N__2731;
    wire N__2726;
    wire N__2723;
    wire N__2720;
    wire N__2719;
    wire N__2716;
    wire N__2713;
    wire N__2708;
    wire N__2707;
    wire N__2704;
    wire N__2701;
    wire N__2696;
    wire N__2695;
    wire N__2692;
    wire N__2689;
    wire N__2686;
    wire N__2681;
    wire N__2680;
    wire N__2677;
    wire N__2674;
    wire N__2669;
    wire N__2668;
    wire N__2665;
    wire N__2662;
    wire N__2657;
    wire N__2656;
    wire N__2653;
    wire N__2650;
    wire N__2645;
    wire N__2644;
    wire N__2641;
    wire N__2638;
    wire N__2635;
    wire N__2630;
    wire N__2629;
    wire N__2626;
    wire N__2623;
    wire N__2618;
    wire N__2615;
    wire N__2612;
    wire N__2609;
    wire N__2606;
    wire N__2603;
    wire N__2602;
    wire N__2599;
    wire N__2596;
    wire N__2591;
    wire N__2588;
    wire N__2585;
    wire N__2582;
    wire N__2579;
    wire N__2576;
    wire N__2573;
    wire N__2570;
    wire N__2567;
    wire N__2566;
    wire N__2563;
    wire N__2560;
    wire N__2557;
    wire N__2552;
    wire N__2549;
    wire N__2546;
    wire N__2543;
    wire N__2540;
    wire N__2537;
    wire N__2534;
    wire N__2531;
    wire N__2528;
    wire N__2525;
    wire N__2522;
    wire N__2521;
    wire N__2520;
    wire N__2519;
    wire N__2518;
    wire N__2515;
    wire N__2512;
    wire N__2509;
    wire N__2504;
    wire N__2495;
    wire N__2492;
    wire N__2491;
    wire N__2488;
    wire N__2485;
    wire N__2480;
    wire N__2479;
    wire N__2476;
    wire N__2475;
    wire N__2474;
    wire N__2471;
    wire N__2470;
    wire N__2467;
    wire N__2464;
    wire N__2461;
    wire N__2456;
    wire N__2447;
    wire N__2444;
    wire N__2443;
    wire N__2440;
    wire N__2437;
    wire N__2432;
    wire N__2431;
    wire N__2430;
    wire N__2429;
    wire N__2428;
    wire N__2425;
    wire N__2422;
    wire N__2419;
    wire N__2414;
    wire N__2405;
    wire N__2404;
    wire N__2403;
    wire N__2396;
    wire N__2393;
    wire N__2390;
    wire N__2389;
    wire N__2386;
    wire N__2383;
    wire N__2378;
    wire N__2377;
    wire N__2376;
    wire N__2373;
    wire N__2372;
    wire N__2371;
    wire N__2368;
    wire N__2365;
    wire N__2362;
    wire N__2359;
    wire N__2356;
    wire N__2345;
    wire N__2342;
    wire N__2339;
    wire N__2336;
    wire N__2333;
    wire N__2332;
    wire N__2329;
    wire N__2326;
    wire N__2323;
    wire N__2318;
    wire N__2317;
    wire N__2314;
    wire N__2311;
    wire N__2306;
    wire N__2303;
    wire N__2302;
    wire N__2297;
    wire N__2294;
    wire N__2291;
    wire N__2288;
    wire N__2285;
    wire N__2284;
    wire N__2281;
    wire N__2278;
    wire N__2275;
    wire N__2272;
    wire N__2267;
    wire N__2264;
    wire N__2263;
    wire N__2260;
    wire N__2257;
    wire N__2254;
    wire N__2249;
    wire N__2246;
    wire N__2243;
    wire N__2240;
    wire N__2237;
    wire N__2234;
    wire N__2231;
    wire N__2228;
    wire N__2227;
    wire N__2224;
    wire N__2223;
    wire N__2220;
    wire N__2217;
    wire N__2214;
    wire N__2213;
    wire N__2210;
    wire N__2205;
    wire N__2202;
    wire N__2195;
    wire N__2192;
    wire N__2189;
    wire N__2186;
    wire N__2185;
    wire N__2180;
    wire N__2177;
    wire N__2176;
    wire N__2171;
    wire N__2168;
    wire N__2165;
    wire N__2164;
    wire N__2159;
    wire N__2156;
    wire N__2155;
    wire N__2150;
    wire N__2147;
    wire N__2144;
    wire N__2141;
    wire N__2138;
    wire N__2135;
    wire N__2132;
    wire N__2129;
    wire N__2126;
    wire N__2123;
    wire N__2120;
    wire N__2117;
    wire N__2114;
    wire N__2111;
    wire N__2108;
    wire N__2105;
    wire N__2102;
    wire N__2099;
    wire N__2096;
    wire N__2093;
    wire N__2090;
    wire N__2087;
    wire N__2084;
    wire N__2081;
    wire N__2078;
    wire N__2075;
    wire N__2072;
    wire N__2069;
    wire N__2066;
    wire N__2065;
    wire N__2060;
    wire N__2057;
    wire N__2056;
    wire N__2053;
    wire N__2050;
    wire N__2045;
    wire N__2042;
    wire N__2041;
    wire N__2038;
    wire N__2033;
    wire N__2030;
    wire N__2029;
    wire N__2026;
    wire N__2021;
    wire N__2018;
    wire N__2017;
    wire N__2014;
    wire N__2009;
    wire N__2006;
    wire N__2003;
    wire N__2002;
    wire N__1999;
    wire N__1996;
    wire N__1991;
    wire N__1990;
    wire N__1987;
    wire N__1984;
    wire N__1979;
    wire N__1976;
    wire N__1975;
    wire N__1970;
    wire N__1967;
    wire N__1966;
    wire N__1963;
    wire N__1958;
    wire N__1955;
    wire N__1954;
    wire N__1949;
    wire N__1946;
    wire N__1945;
    wire N__1940;
    wire N__1937;
    wire N__1936;
    wire N__1931;
    wire N__1928;
    wire N__1925;
    wire N__1924;
    wire N__1919;
    wire N__1916;
    wire N__1915;
    wire N__1910;
    wire N__1907;
    wire N__1906;
    wire N__1903;
    wire N__1900;
    wire N__1897;
    wire N__1892;
    wire N__1889;
    wire N__1886;
    wire N__1883;
    wire N__1880;
    wire N__1879;
    wire N__1876;
    wire N__1873;
    wire N__1872;
    wire N__1869;
    wire N__1866;
    wire N__1863;
    wire N__1856;
    wire N__1853;
    wire N__1850;
    wire N__1847;
    wire N__1844;
    wire N__1841;
    wire io_jtag_tck_pad_gb_input;
    wire VCCG0;
    wire GNDG0;
    wire io_leds_c_0;
    wire ctrl_idcodeArea_shifter_7;
    wire ctrl_idcodeArea_shifter_10;
    wire ctrl_idcodeArea_shifter_9;
    wire ctrl_idcodeArea_shifter_8;
    wire ctrl_idcodeArea_shifter_4;
    wire ctrl_idcodeArea_shifter_6;
    wire ctrl_idcodeArea_shifter_5;
    wire ctrl_idcodeArea_shifter_11;
    wire ctrl_idcodeArea_shifter_16;
    wire ctrl_idcodeArea_shifter_15;
    wire ctrl_idcodeArea_shifter_14;
    wire ctrl_idcodeArea_shifter_13;
    wire ctrl_idcodeArea_shifter_12;
    wire ctrl_idcodeArea_shifter_3;
    wire ctrl_idcodeArea_shifter_2;
    wire n7;
    wire n7_cascade_;
    wire n2206;
    wire n7_adj_1_cascade_;
    wire bfn_4_7_0_;
    wire n2059;
    wire n2060;
    wire n2061;
    wire n2062;
    wire n2063;
    wire n2064;
    wire n2065;
    wire n2066;
    wire bfn_4_8_0_;
    wire n2067;
    wire n2068;
    wire n2069;
    wire n2070;
    wire n2071;
    wire n2072;
    wire n2073;
    wire n2074;
    wire bfn_4_9_0_;
    wire n2075;
    wire n2076;
    wire n2077;
    wire n2078;
    wire n2079;
    wire n2080;
    wire global_reset_c;
    wire ctrl_idcodeArea_shifter_31;
    wire ctrl_idcodeArea_shifter_28;
    wire ctrl_idcodeArea_shifter_30;
    wire ctrl_idcodeArea_shifter_29;
    wire ctrl_idcodeArea_shifter_17;
    wire ctrl_idcodeArea_shifter_1;
    wire n6_cascade_;
    wire ctrl_idcodeArea_shifter_0;
    wire n2085;
    wire n15_cascade_;
    wire n7_adj_1;
    wire ctrl_ledsArea_shifter_0;
    wire ctrl_tap_tdoUnbufferd_N_211_cascade_;
    wire ctrl_tap_tdoUnbufferd;
    wire n1489_cascade_;
    wire n1269_cascade_;
    wire ctrl_tap_instruction_0;
    wire ctrl_tap_instructionShift_3;
    wire ctrl_tap_instruction_3;
    wire ctrl_tap_instructionShift_2;
    wire ctrl_tap_instruction_2;
    wire n1269;
    wire ctrl_tap_instructionShift_1;
    wire ctrl_tap_instruction_1;
    wire n2248;
    wire n118_cascade_;
    wire n2282_cascade_;
    wire n2326_cascade_;
    wire n2306;
    wire n1022;
    wire n2231_cascade_;
    wire n2273;
    wire n2263_cascade_;
    wire n2323;
    wire n2272;
    wire io_leds_c_7;
    wire myClockArea_timeout_counter_value_3;
    wire myClockArea_timeout_counter_value_1;
    wire myClockArea_timeout_counter_value_5;
    wire myClockArea_timeout_counter_value_0;
    wire n2309;
    wire myClockArea_timeout_counter_value_4;
    wire myClockArea_timeout_counter_value_6;
    wire myClockArea_timeout_counter_value_22;
    wire myClockArea_timeout_counter_value_16;
    wire myClockArea_timeout_counter_value_17;
    wire myClockArea_timeout_counter_value_8;
    wire myClockArea_timeout_counter_value_10;
    wire myClockArea_timeout_counter_value_2;
    wire n2216;
    wire n2218_cascade_;
    wire n2222;
    wire myClockArea_timeout_counter_value_13;
    wire n2228_cascade_;
    wire n2185;
    wire n2185_cascade_;
    wire n1848;
    wire myClockArea_timeout_counter_value_7;
    wire myClockArea_timeout_counter_value_21;
    wire n11;
    wire myClockArea_timeout_counter_value_19;
    wire myClockArea_timeout_counter_value_15;
    wire myClockArea_timeout_counter_value_20;
    wire myClockArea_timeout_counter_value_11;
    wire n2220;
    wire myClockArea_timeout_counter_value_9;
    wire myClockArea_timeout_counter_value_18;
    wire myClockArea_timeout_counter_value_12;
    wire myClockArea_timeout_counter_value_14;
    wire n13;
    wire myClockArea_timeout_state;
    wire io_leds_c_3;
    wire global_clk_c;
    wire ctrl_idcodeArea_shifter_25;
    wire ctrl_idcodeArea_shifter_24;
    wire ctrl_idcodeArea_shifter_27;
    wire ctrl_idcodeArea_shifter_26;
    wire io_jtag_tdi_c;
    wire ctrl_idcodeArea_shifter_23;
    wire ctrl_idcodeArea_shifter_22;
    wire ctrl_idcodeArea_shifter_21;
    wire ctrl_idcodeArea_shifter_18;
    wire n15;
    wire ctrl_idcodeArea_shifter_20;
    wire n1489;
    wire ctrl_idcodeArea_shifter_19;
    wire n17_cascade_;
    wire n1687_cascade_;
    wire n2234;
    wire n8;
    wire n2198;
    wire ctrl_tap_instructionShift_0;
    wire ctrl_tap_bypass;
    wire n2198_cascade_;
    wire n4;
    wire ctrl_tap_tdoUnbufferd_N_213;
    wire n1686;
    wire n112_cascade_;
    wire n929;
    wire n1117;
    wire n2260_cascade_;
    wire n1119;
    wire ctrl_tap_fsm_state_3;
    wire ctrl_tap_fsm_state_2;
    wire ctrl_tap_fsm_stateNext_3__N_10_c_3;
    wire ctrl_tap_fsm_state_1;
    wire n2243;
    wire n2186;
    wire ctrl_tap_fsm_state_0;
    wire io_leds_c_1;
    wire ctrl_ledsArea_shifter_1;
    wire ctrl_ledsArea_store_3;
    wire ctrl_ledsArea_shifter_3;
    wire io_leds_c_5;
    wire ctrl_ledsArea_shifter_5;
    wire ctrl_ledsArea_shifter_7;
    wire n1638;
    wire io_leds_c_6;
    wire n7_adj_2;
    wire ctrl_ledsArea_shifter_6;
    wire n1275;
    wire ctrl_ledsArea_shifter_4;
    wire io_leds_c_4;
    wire ctrl_ledsArea_shifter_2;
    wire n2110;
    wire io_leds_c_2;
    wire io_jtag_tck_c;
    wire _gnd_net_;

    PRE_IO_GBUF global_clk_pad_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__4908),
            .GLOBALBUFFEROUTPUT(global_clk_c));
    defparam global_clk_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam global_clk_pad_iopad.PULLUP=1'b0;
    IO_PAD global_clk_pad_iopad (
            .OE(N__4910),
            .DIN(N__4909),
            .DOUT(N__4908),
            .PACKAGEPIN(global_clk));
    defparam global_clk_pad_preio.PIN_TYPE=6'b000001;
    defparam global_clk_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO global_clk_pad_preio (
            .PADOEN(N__4910),
            .PADOUT(N__4909),
            .PADIN(N__4908),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam ctrl_tap_fsm_stateNext_3__N_10_pad_3_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ctrl_tap_fsm_stateNext_3__N_10_pad_3_iopad.PULLUP=1'b0;
    IO_PAD ctrl_tap_fsm_stateNext_3__N_10_pad_3_iopad (
            .OE(N__4899),
            .DIN(N__4898),
            .DOUT(N__4897),
            .PACKAGEPIN(io_jtag_tms));
    defparam ctrl_tap_fsm_stateNext_3__N_10_pad_3_preio.PIN_TYPE=6'b000001;
    defparam ctrl_tap_fsm_stateNext_3__N_10_pad_3_preio.NEG_TRIGGER=1'b0;
    PRE_IO ctrl_tap_fsm_stateNext_3__N_10_pad_3_preio (
            .PADOEN(N__4899),
            .PADOUT(N__4898),
            .PADIN(N__4897),
            .CLOCKENABLE(),
            .DIN0(ctrl_tap_fsm_stateNext_3__N_10_c_3),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam global_reset_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam global_reset_pad_iopad.PULLUP=1'b0;
    IO_PAD global_reset_pad_iopad (
            .OE(N__4890),
            .DIN(N__4889),
            .DOUT(N__4888),
            .PACKAGEPIN(global_reset));
    defparam global_reset_pad_preio.PIN_TYPE=6'b000001;
    defparam global_reset_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO global_reset_pad_preio (
            .PADOEN(N__4890),
            .PADOUT(N__4889),
            .PADIN(N__4888),
            .CLOCKENABLE(),
            .DIN0(global_reset_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam io_jtag_tdi_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam io_jtag_tdi_pad_iopad.PULLUP=1'b0;
    IO_PAD io_jtag_tdi_pad_iopad (
            .OE(N__4881),
            .DIN(N__4880),
            .DOUT(N__4879),
            .PACKAGEPIN(io_jtag_tdi));
    defparam io_jtag_tdi_pad_preio.PIN_TYPE=6'b000001;
    defparam io_jtag_tdi_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO io_jtag_tdi_pad_preio (
            .PADOEN(N__4881),
            .PADOUT(N__4880),
            .PADIN(N__4879),
            .CLOCKENABLE(),
            .DIN0(io_jtag_tdi_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam io_jtag_tdo_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam io_jtag_tdo_pad_iopad.PULLUP=1'b0;
    IO_PAD io_jtag_tdo_pad_iopad (
            .OE(N__4872),
            .DIN(N__4871),
            .DOUT(N__4870),
            .PACKAGEPIN(io_jtag_tdo));
    defparam io_jtag_tdo_pad_preio.PIN_TYPE=6'b010101;
    defparam io_jtag_tdo_pad_preio.NEG_TRIGGER=1'b1;
    PRE_IO io_jtag_tdo_pad_preio (
            .PADOEN(N__4872),
            .PADOUT(N__4871),
            .PADIN(N__4870),
            .CLOCKENABLE(VCCG0),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__2246),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(N__4322),
            .OUTPUTENABLE());
    defparam io_leds_pad_0_iopad.IO_STANDARD="SB_LVCMOS";
    defparam io_leds_pad_0_iopad.PULLUP=1'b0;
    IO_PAD io_leds_pad_0_iopad (
            .OE(N__4863),
            .DIN(N__4862),
            .DOUT(N__4861),
            .PACKAGEPIN(io_leds[0]));
    defparam io_leds_pad_0_preio.PIN_TYPE=6'b011001;
    defparam io_leds_pad_0_preio.NEG_TRIGGER=1'b0;
    PRE_IO io_leds_pad_0_preio (
            .PADOEN(N__4863),
            .PADOUT(N__4862),
            .PADIN(N__4861),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__1892),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam io_leds_pad_1_iopad.IO_STANDARD="SB_LVCMOS";
    defparam io_leds_pad_1_iopad.PULLUP=1'b0;
    IO_PAD io_leds_pad_1_iopad (
            .OE(N__4854),
            .DIN(N__4853),
            .DOUT(N__4852),
            .PACKAGEPIN(io_leds[1]));
    defparam io_leds_pad_1_preio.PIN_TYPE=6'b011001;
    defparam io_leds_pad_1_preio.NEG_TRIGGER=1'b0;
    PRE_IO io_leds_pad_1_preio (
            .PADOEN(N__4854),
            .PADOUT(N__4853),
            .PADIN(N__4852),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__4772),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam io_leds_pad_2_iopad.IO_STANDARD="SB_LVCMOS";
    defparam io_leds_pad_2_iopad.PULLUP=1'b0;
    IO_PAD io_leds_pad_2_iopad (
            .OE(N__4845),
            .DIN(N__4844),
            .DOUT(N__4843),
            .PACKAGEPIN(io_leds[2]));
    defparam io_leds_pad_2_preio.PIN_TYPE=6'b011001;
    defparam io_leds_pad_2_preio.NEG_TRIGGER=1'b0;
    PRE_IO io_leds_pad_2_preio (
            .PADOEN(N__4845),
            .PADOUT(N__4844),
            .PADIN(N__4843),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__4355),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam io_leds_pad_3_iopad.IO_STANDARD="SB_LVCMOS";
    defparam io_leds_pad_3_iopad.PULLUP=1'b0;
    IO_PAD io_leds_pad_3_iopad (
            .OE(N__4836),
            .DIN(N__4835),
            .DOUT(N__4834),
            .PACKAGEPIN(io_leds[3]));
    defparam io_leds_pad_3_preio.PIN_TYPE=6'b011001;
    defparam io_leds_pad_3_preio.NEG_TRIGGER=1'b0;
    PRE_IO io_leds_pad_3_preio (
            .PADOEN(N__4836),
            .PADOUT(N__4835),
            .PADIN(N__4834),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__2864),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam io_leds_pad_4_iopad.IO_STANDARD="SB_LVCMOS";
    defparam io_leds_pad_4_iopad.PULLUP=1'b0;
    IO_PAD io_leds_pad_4_iopad (
            .OE(N__4827),
            .DIN(N__4826),
            .DOUT(N__4825),
            .PACKAGEPIN(io_leds[4]));
    defparam io_leds_pad_4_preio.PIN_TYPE=6'b011001;
    defparam io_leds_pad_4_preio.NEG_TRIGGER=1'b0;
    PRE_IO io_leds_pad_4_preio (
            .PADOEN(N__4827),
            .PADOUT(N__4826),
            .PADIN(N__4825),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__4457),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam io_leds_pad_5_iopad.IO_STANDARD="SB_LVCMOS";
    defparam io_leds_pad_5_iopad.PULLUP=1'b0;
    IO_PAD io_leds_pad_5_iopad (
            .OE(N__4818),
            .DIN(N__4817),
            .DOUT(N__4816),
            .PACKAGEPIN(io_leds[5]));
    defparam io_leds_pad_5_preio.PIN_TYPE=6'b011001;
    defparam io_leds_pad_5_preio.NEG_TRIGGER=1'b0;
    PRE_IO io_leds_pad_5_preio (
            .PADOEN(N__4818),
            .PADOUT(N__4817),
            .PADIN(N__4816),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__4697),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam io_leds_pad_6_iopad.IO_STANDARD="SB_LVCMOS";
    defparam io_leds_pad_6_iopad.PULLUP=1'b0;
    IO_PAD io_leds_pad_6_iopad (
            .OE(N__4809),
            .DIN(N__4808),
            .DOUT(N__4807),
            .PACKAGEPIN(io_leds[6]));
    defparam io_leds_pad_6_preio.PIN_TYPE=6'b011001;
    defparam io_leds_pad_6_preio.NEG_TRIGGER=1'b0;
    PRE_IO io_leds_pad_6_preio (
            .PADOEN(N__4809),
            .PADOUT(N__4808),
            .PADIN(N__4807),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__4607),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam io_leds_pad_7_iopad.IO_STANDARD="SB_LVCMOS";
    defparam io_leds_pad_7_iopad.PULLUP=1'b0;
    IO_PAD io_leds_pad_7_iopad (
            .OE(N__4800),
            .DIN(N__4799),
            .DOUT(N__4798),
            .PACKAGEPIN(io_leds[7]));
    defparam io_leds_pad_7_preio.PIN_TYPE=6'b011001;
    defparam io_leds_pad_7_preio.NEG_TRIGGER=1'b0;
    PRE_IO io_leds_pad_7_preio (
            .PADOEN(N__4800),
            .PADOUT(N__4799),
            .PADIN(N__4798),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__2807),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam io_jtag_tck_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam io_jtag_tck_pad_iopad.PULLUP=1'b0;
    IO_PAD io_jtag_tck_pad_iopad (
            .OE(N__4791),
            .DIN(N__4790),
            .DOUT(N__4789),
            .PACKAGEPIN(io_jtag_tck));
    defparam io_jtag_tck_pad_preio.PIN_TYPE=6'b000001;
    defparam io_jtag_tck_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO io_jtag_tck_pad_preio (
            .PADOEN(N__4791),
            .PADOUT(N__4790),
            .PADIN(N__4789),
            .CLOCKENABLE(),
            .DIN0(io_jtag_tck_pad_gb_input),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IoInMux I__1134 (
            .O(N__4772),
            .I(N__4769));
    LocalMux I__1133 (
            .O(N__4769),
            .I(N__4766));
    IoSpan4Mux I__1132 (
            .O(N__4766),
            .I(N__4763));
    Span4Mux_s2_h I__1131 (
            .O(N__4763),
            .I(N__4759));
    CascadeMux I__1130 (
            .O(N__4762),
            .I(N__4756));
    Span4Mux_h I__1129 (
            .O(N__4759),
            .I(N__4752));
    InMux I__1128 (
            .O(N__4756),
            .I(N__4749));
    InMux I__1127 (
            .O(N__4755),
            .I(N__4746));
    Odrv4 I__1126 (
            .O(N__4752),
            .I(io_leds_c_1));
    LocalMux I__1125 (
            .O(N__4749),
            .I(io_leds_c_1));
    LocalMux I__1124 (
            .O(N__4746),
            .I(io_leds_c_1));
    InMux I__1123 (
            .O(N__4739),
            .I(N__4735));
    InMux I__1122 (
            .O(N__4738),
            .I(N__4732));
    LocalMux I__1121 (
            .O(N__4735),
            .I(N__4729));
    LocalMux I__1120 (
            .O(N__4732),
            .I(ctrl_ledsArea_shifter_1));
    Odrv12 I__1119 (
            .O(N__4729),
            .I(ctrl_ledsArea_shifter_1));
    CascadeMux I__1118 (
            .O(N__4724),
            .I(N__4721));
    InMux I__1117 (
            .O(N__4721),
            .I(N__4717));
    InMux I__1116 (
            .O(N__4720),
            .I(N__4714));
    LocalMux I__1115 (
            .O(N__4717),
            .I(ctrl_ledsArea_store_3));
    LocalMux I__1114 (
            .O(N__4714),
            .I(ctrl_ledsArea_store_3));
    InMux I__1113 (
            .O(N__4709),
            .I(N__4705));
    InMux I__1112 (
            .O(N__4708),
            .I(N__4702));
    LocalMux I__1111 (
            .O(N__4705),
            .I(ctrl_ledsArea_shifter_3));
    LocalMux I__1110 (
            .O(N__4702),
            .I(ctrl_ledsArea_shifter_3));
    IoInMux I__1109 (
            .O(N__4697),
            .I(N__4693));
    CascadeMux I__1108 (
            .O(N__4696),
            .I(N__4690));
    LocalMux I__1107 (
            .O(N__4693),
            .I(N__4687));
    InMux I__1106 (
            .O(N__4690),
            .I(N__4684));
    IoSpan4Mux I__1105 (
            .O(N__4687),
            .I(N__4681));
    LocalMux I__1104 (
            .O(N__4684),
            .I(N__4678));
    Span4Mux_s3_h I__1103 (
            .O(N__4681),
            .I(N__4672));
    Span4Mux_v I__1102 (
            .O(N__4678),
            .I(N__4672));
    InMux I__1101 (
            .O(N__4677),
            .I(N__4669));
    Odrv4 I__1100 (
            .O(N__4672),
            .I(io_leds_c_5));
    LocalMux I__1099 (
            .O(N__4669),
            .I(io_leds_c_5));
    InMux I__1098 (
            .O(N__4664),
            .I(N__4660));
    CascadeMux I__1097 (
            .O(N__4663),
            .I(N__4657));
    LocalMux I__1096 (
            .O(N__4660),
            .I(N__4654));
    InMux I__1095 (
            .O(N__4657),
            .I(N__4651));
    Span4Mux_h I__1094 (
            .O(N__4654),
            .I(N__4648));
    LocalMux I__1093 (
            .O(N__4651),
            .I(ctrl_ledsArea_shifter_5));
    Odrv4 I__1092 (
            .O(N__4648),
            .I(ctrl_ledsArea_shifter_5));
    InMux I__1091 (
            .O(N__4643),
            .I(N__4639));
    InMux I__1090 (
            .O(N__4642),
            .I(N__4636));
    LocalMux I__1089 (
            .O(N__4639),
            .I(N__4633));
    LocalMux I__1088 (
            .O(N__4636),
            .I(ctrl_ledsArea_shifter_7));
    Odrv12 I__1087 (
            .O(N__4633),
            .I(ctrl_ledsArea_shifter_7));
    InMux I__1086 (
            .O(N__4628),
            .I(N__4619));
    InMux I__1085 (
            .O(N__4627),
            .I(N__4619));
    InMux I__1084 (
            .O(N__4626),
            .I(N__4612));
    InMux I__1083 (
            .O(N__4625),
            .I(N__4612));
    InMux I__1082 (
            .O(N__4624),
            .I(N__4612));
    LocalMux I__1081 (
            .O(N__4619),
            .I(n1638));
    LocalMux I__1080 (
            .O(N__4612),
            .I(n1638));
    IoInMux I__1079 (
            .O(N__4607),
            .I(N__4604));
    LocalMux I__1078 (
            .O(N__4604),
            .I(N__4601));
    IoSpan4Mux I__1077 (
            .O(N__4601),
            .I(N__4597));
    CascadeMux I__1076 (
            .O(N__4600),
            .I(N__4594));
    Span4Mux_s0_h I__1075 (
            .O(N__4597),
            .I(N__4591));
    InMux I__1074 (
            .O(N__4594),
            .I(N__4588));
    Span4Mux_h I__1073 (
            .O(N__4591),
            .I(N__4583));
    LocalMux I__1072 (
            .O(N__4588),
            .I(N__4583));
    Span4Mux_h I__1071 (
            .O(N__4583),
            .I(N__4579));
    InMux I__1070 (
            .O(N__4582),
            .I(N__4576));
    Odrv4 I__1069 (
            .O(N__4579),
            .I(io_leds_c_6));
    LocalMux I__1068 (
            .O(N__4576),
            .I(io_leds_c_6));
    InMux I__1067 (
            .O(N__4571),
            .I(N__4567));
    InMux I__1066 (
            .O(N__4570),
            .I(N__4564));
    LocalMux I__1065 (
            .O(N__4567),
            .I(N__4561));
    LocalMux I__1064 (
            .O(N__4564),
            .I(N__4558));
    Span4Mux_v I__1063 (
            .O(N__4561),
            .I(N__4548));
    Span4Mux_v I__1062 (
            .O(N__4558),
            .I(N__4545));
    InMux I__1061 (
            .O(N__4557),
            .I(N__4534));
    InMux I__1060 (
            .O(N__4556),
            .I(N__4534));
    InMux I__1059 (
            .O(N__4555),
            .I(N__4534));
    InMux I__1058 (
            .O(N__4554),
            .I(N__4534));
    InMux I__1057 (
            .O(N__4553),
            .I(N__4534));
    InMux I__1056 (
            .O(N__4552),
            .I(N__4529));
    InMux I__1055 (
            .O(N__4551),
            .I(N__4529));
    Odrv4 I__1054 (
            .O(N__4548),
            .I(n7_adj_2));
    Odrv4 I__1053 (
            .O(N__4545),
            .I(n7_adj_2));
    LocalMux I__1052 (
            .O(N__4534),
            .I(n7_adj_2));
    LocalMux I__1051 (
            .O(N__4529),
            .I(n7_adj_2));
    InMux I__1050 (
            .O(N__4520),
            .I(N__4517));
    LocalMux I__1049 (
            .O(N__4517),
            .I(N__4514));
    Span4Mux_h I__1048 (
            .O(N__4514),
            .I(N__4510));
    InMux I__1047 (
            .O(N__4513),
            .I(N__4507));
    Odrv4 I__1046 (
            .O(N__4510),
            .I(ctrl_ledsArea_shifter_6));
    LocalMux I__1045 (
            .O(N__4507),
            .I(ctrl_ledsArea_shifter_6));
    CEMux I__1044 (
            .O(N__4502),
            .I(N__4499));
    LocalMux I__1043 (
            .O(N__4499),
            .I(N__4494));
    CEMux I__1042 (
            .O(N__4498),
            .I(N__4491));
    CEMux I__1041 (
            .O(N__4497),
            .I(N__4488));
    Span4Mux_h I__1040 (
            .O(N__4494),
            .I(N__4485));
    LocalMux I__1039 (
            .O(N__4491),
            .I(N__4482));
    LocalMux I__1038 (
            .O(N__4488),
            .I(N__4479));
    Odrv4 I__1037 (
            .O(N__4485),
            .I(n1275));
    Odrv4 I__1036 (
            .O(N__4482),
            .I(n1275));
    Odrv4 I__1035 (
            .O(N__4479),
            .I(n1275));
    InMux I__1034 (
            .O(N__4472),
            .I(N__4468));
    InMux I__1033 (
            .O(N__4471),
            .I(N__4465));
    LocalMux I__1032 (
            .O(N__4468),
            .I(N__4462));
    LocalMux I__1031 (
            .O(N__4465),
            .I(ctrl_ledsArea_shifter_4));
    Odrv4 I__1030 (
            .O(N__4462),
            .I(ctrl_ledsArea_shifter_4));
    IoInMux I__1029 (
            .O(N__4457),
            .I(N__4454));
    LocalMux I__1028 (
            .O(N__4454),
            .I(N__4451));
    Span12Mux_s5_h I__1027 (
            .O(N__4451),
            .I(N__4446));
    InMux I__1026 (
            .O(N__4450),
            .I(N__4443));
    InMux I__1025 (
            .O(N__4449),
            .I(N__4440));
    Odrv12 I__1024 (
            .O(N__4446),
            .I(io_leds_c_4));
    LocalMux I__1023 (
            .O(N__4443),
            .I(io_leds_c_4));
    LocalMux I__1022 (
            .O(N__4440),
            .I(io_leds_c_4));
    InMux I__1021 (
            .O(N__4433),
            .I(N__4430));
    LocalMux I__1020 (
            .O(N__4430),
            .I(N__4426));
    InMux I__1019 (
            .O(N__4429),
            .I(N__4423));
    Odrv4 I__1018 (
            .O(N__4426),
            .I(ctrl_ledsArea_shifter_2));
    LocalMux I__1017 (
            .O(N__4423),
            .I(ctrl_ledsArea_shifter_2));
    InMux I__1016 (
            .O(N__4418),
            .I(N__4411));
    InMux I__1015 (
            .O(N__4417),
            .I(N__4408));
    InMux I__1014 (
            .O(N__4416),
            .I(N__4405));
    InMux I__1013 (
            .O(N__4415),
            .I(N__4402));
    InMux I__1012 (
            .O(N__4414),
            .I(N__4397));
    LocalMux I__1011 (
            .O(N__4411),
            .I(N__4394));
    LocalMux I__1010 (
            .O(N__4408),
            .I(N__4388));
    LocalMux I__1009 (
            .O(N__4405),
            .I(N__4388));
    LocalMux I__1008 (
            .O(N__4402),
            .I(N__4385));
    InMux I__1007 (
            .O(N__4401),
            .I(N__4380));
    InMux I__1006 (
            .O(N__4400),
            .I(N__4380));
    LocalMux I__1005 (
            .O(N__4397),
            .I(N__4377));
    Span4Mux_h I__1004 (
            .O(N__4394),
            .I(N__4374));
    InMux I__1003 (
            .O(N__4393),
            .I(N__4371));
    Span4Mux_v I__1002 (
            .O(N__4388),
            .I(N__4364));
    Span4Mux_v I__1001 (
            .O(N__4385),
            .I(N__4364));
    LocalMux I__1000 (
            .O(N__4380),
            .I(N__4364));
    Odrv4 I__999 (
            .O(N__4377),
            .I(n2110));
    Odrv4 I__998 (
            .O(N__4374),
            .I(n2110));
    LocalMux I__997 (
            .O(N__4371),
            .I(n2110));
    Odrv4 I__996 (
            .O(N__4364),
            .I(n2110));
    IoInMux I__995 (
            .O(N__4355),
            .I(N__4352));
    LocalMux I__994 (
            .O(N__4352),
            .I(N__4348));
    CascadeMux I__993 (
            .O(N__4351),
            .I(N__4345));
    IoSpan4Mux I__992 (
            .O(N__4348),
            .I(N__4342));
    InMux I__991 (
            .O(N__4345),
            .I(N__4339));
    Span4Mux_s2_h I__990 (
            .O(N__4342),
            .I(N__4335));
    LocalMux I__989 (
            .O(N__4339),
            .I(N__4332));
    InMux I__988 (
            .O(N__4338),
            .I(N__4329));
    Odrv4 I__987 (
            .O(N__4335),
            .I(io_leds_c_2));
    Odrv4 I__986 (
            .O(N__4332),
            .I(io_leds_c_2));
    LocalMux I__985 (
            .O(N__4329),
            .I(io_leds_c_2));
    ClkMux I__984 (
            .O(N__4322),
            .I(N__4265));
    ClkMux I__983 (
            .O(N__4321),
            .I(N__4265));
    ClkMux I__982 (
            .O(N__4320),
            .I(N__4265));
    ClkMux I__981 (
            .O(N__4319),
            .I(N__4265));
    ClkMux I__980 (
            .O(N__4318),
            .I(N__4265));
    ClkMux I__979 (
            .O(N__4317),
            .I(N__4265));
    ClkMux I__978 (
            .O(N__4316),
            .I(N__4265));
    ClkMux I__977 (
            .O(N__4315),
            .I(N__4265));
    ClkMux I__976 (
            .O(N__4314),
            .I(N__4265));
    ClkMux I__975 (
            .O(N__4313),
            .I(N__4265));
    ClkMux I__974 (
            .O(N__4312),
            .I(N__4265));
    ClkMux I__973 (
            .O(N__4311),
            .I(N__4265));
    ClkMux I__972 (
            .O(N__4310),
            .I(N__4265));
    ClkMux I__971 (
            .O(N__4309),
            .I(N__4265));
    ClkMux I__970 (
            .O(N__4308),
            .I(N__4265));
    ClkMux I__969 (
            .O(N__4307),
            .I(N__4265));
    ClkMux I__968 (
            .O(N__4306),
            .I(N__4265));
    ClkMux I__967 (
            .O(N__4305),
            .I(N__4265));
    ClkMux I__966 (
            .O(N__4304),
            .I(N__4265));
    GlobalMux I__965 (
            .O(N__4265),
            .I(N__4262));
    gio2CtrlBuf I__964 (
            .O(N__4262),
            .I(io_jtag_tck_c));
    InMux I__963 (
            .O(N__4259),
            .I(N__4255));
    InMux I__962 (
            .O(N__4258),
            .I(N__4252));
    LocalMux I__961 (
            .O(N__4255),
            .I(n1686));
    LocalMux I__960 (
            .O(N__4252),
            .I(n1686));
    CascadeMux I__959 (
            .O(N__4247),
            .I(n112_cascade_));
    InMux I__958 (
            .O(N__4244),
            .I(N__4241));
    LocalMux I__957 (
            .O(N__4241),
            .I(N__4238));
    Odrv4 I__956 (
            .O(N__4238),
            .I(n929));
    CascadeMux I__955 (
            .O(N__4235),
            .I(N__4232));
    InMux I__954 (
            .O(N__4232),
            .I(N__4228));
    InMux I__953 (
            .O(N__4231),
            .I(N__4223));
    LocalMux I__952 (
            .O(N__4228),
            .I(N__4220));
    InMux I__951 (
            .O(N__4227),
            .I(N__4215));
    InMux I__950 (
            .O(N__4226),
            .I(N__4215));
    LocalMux I__949 (
            .O(N__4223),
            .I(n1117));
    Odrv4 I__948 (
            .O(N__4220),
            .I(n1117));
    LocalMux I__947 (
            .O(N__4215),
            .I(n1117));
    CascadeMux I__946 (
            .O(N__4208),
            .I(n2260_cascade_));
    InMux I__945 (
            .O(N__4205),
            .I(N__4195));
    InMux I__944 (
            .O(N__4204),
            .I(N__4192));
    InMux I__943 (
            .O(N__4203),
            .I(N__4189));
    InMux I__942 (
            .O(N__4202),
            .I(N__4184));
    InMux I__941 (
            .O(N__4201),
            .I(N__4184));
    InMux I__940 (
            .O(N__4200),
            .I(N__4181));
    InMux I__939 (
            .O(N__4199),
            .I(N__4178));
    InMux I__938 (
            .O(N__4198),
            .I(N__4175));
    LocalMux I__937 (
            .O(N__4195),
            .I(n1119));
    LocalMux I__936 (
            .O(N__4192),
            .I(n1119));
    LocalMux I__935 (
            .O(N__4189),
            .I(n1119));
    LocalMux I__934 (
            .O(N__4184),
            .I(n1119));
    LocalMux I__933 (
            .O(N__4181),
            .I(n1119));
    LocalMux I__932 (
            .O(N__4178),
            .I(n1119));
    LocalMux I__931 (
            .O(N__4175),
            .I(n1119));
    CascadeMux I__930 (
            .O(N__4160),
            .I(N__4157));
    InMux I__929 (
            .O(N__4157),
            .I(N__4145));
    InMux I__928 (
            .O(N__4156),
            .I(N__4145));
    InMux I__927 (
            .O(N__4155),
            .I(N__4145));
    CascadeMux I__926 (
            .O(N__4154),
            .I(N__4137));
    InMux I__925 (
            .O(N__4153),
            .I(N__4134));
    InMux I__924 (
            .O(N__4152),
            .I(N__4131));
    LocalMux I__923 (
            .O(N__4145),
            .I(N__4128));
    CascadeMux I__922 (
            .O(N__4144),
            .I(N__4125));
    CascadeMux I__921 (
            .O(N__4143),
            .I(N__4117));
    InMux I__920 (
            .O(N__4142),
            .I(N__4107));
    InMux I__919 (
            .O(N__4141),
            .I(N__4100));
    InMux I__918 (
            .O(N__4140),
            .I(N__4100));
    InMux I__917 (
            .O(N__4137),
            .I(N__4100));
    LocalMux I__916 (
            .O(N__4134),
            .I(N__4095));
    LocalMux I__915 (
            .O(N__4131),
            .I(N__4095));
    Span4Mux_v I__914 (
            .O(N__4128),
            .I(N__4092));
    InMux I__913 (
            .O(N__4125),
            .I(N__4083));
    InMux I__912 (
            .O(N__4124),
            .I(N__4083));
    InMux I__911 (
            .O(N__4123),
            .I(N__4083));
    InMux I__910 (
            .O(N__4122),
            .I(N__4083));
    InMux I__909 (
            .O(N__4121),
            .I(N__4076));
    InMux I__908 (
            .O(N__4120),
            .I(N__4076));
    InMux I__907 (
            .O(N__4117),
            .I(N__4076));
    InMux I__906 (
            .O(N__4116),
            .I(N__4067));
    InMux I__905 (
            .O(N__4115),
            .I(N__4067));
    InMux I__904 (
            .O(N__4114),
            .I(N__4067));
    InMux I__903 (
            .O(N__4113),
            .I(N__4067));
    InMux I__902 (
            .O(N__4112),
            .I(N__4060));
    InMux I__901 (
            .O(N__4111),
            .I(N__4060));
    InMux I__900 (
            .O(N__4110),
            .I(N__4060));
    LocalMux I__899 (
            .O(N__4107),
            .I(ctrl_tap_fsm_state_3));
    LocalMux I__898 (
            .O(N__4100),
            .I(ctrl_tap_fsm_state_3));
    Odrv4 I__897 (
            .O(N__4095),
            .I(ctrl_tap_fsm_state_3));
    Odrv4 I__896 (
            .O(N__4092),
            .I(ctrl_tap_fsm_state_3));
    LocalMux I__895 (
            .O(N__4083),
            .I(ctrl_tap_fsm_state_3));
    LocalMux I__894 (
            .O(N__4076),
            .I(ctrl_tap_fsm_state_3));
    LocalMux I__893 (
            .O(N__4067),
            .I(ctrl_tap_fsm_state_3));
    LocalMux I__892 (
            .O(N__4060),
            .I(ctrl_tap_fsm_state_3));
    CascadeMux I__891 (
            .O(N__4043),
            .I(N__4029));
    CascadeMux I__890 (
            .O(N__4042),
            .I(N__4024));
    CascadeMux I__889 (
            .O(N__4041),
            .I(N__4018));
    InMux I__888 (
            .O(N__4040),
            .I(N__4010));
    InMux I__887 (
            .O(N__4039),
            .I(N__4010));
    InMux I__886 (
            .O(N__4038),
            .I(N__4010));
    InMux I__885 (
            .O(N__4037),
            .I(N__4007));
    InMux I__884 (
            .O(N__4036),
            .I(N__4004));
    InMux I__883 (
            .O(N__4035),
            .I(N__4001));
    InMux I__882 (
            .O(N__4034),
            .I(N__3996));
    InMux I__881 (
            .O(N__4033),
            .I(N__3996));
    InMux I__880 (
            .O(N__4032),
            .I(N__3987));
    InMux I__879 (
            .O(N__4029),
            .I(N__3987));
    InMux I__878 (
            .O(N__4028),
            .I(N__3987));
    InMux I__877 (
            .O(N__4027),
            .I(N__3987));
    InMux I__876 (
            .O(N__4024),
            .I(N__3980));
    InMux I__875 (
            .O(N__4023),
            .I(N__3980));
    InMux I__874 (
            .O(N__4022),
            .I(N__3980));
    InMux I__873 (
            .O(N__4021),
            .I(N__3973));
    InMux I__872 (
            .O(N__4018),
            .I(N__3973));
    InMux I__871 (
            .O(N__4017),
            .I(N__3973));
    LocalMux I__870 (
            .O(N__4010),
            .I(ctrl_tap_fsm_state_2));
    LocalMux I__869 (
            .O(N__4007),
            .I(ctrl_tap_fsm_state_2));
    LocalMux I__868 (
            .O(N__4004),
            .I(ctrl_tap_fsm_state_2));
    LocalMux I__867 (
            .O(N__4001),
            .I(ctrl_tap_fsm_state_2));
    LocalMux I__866 (
            .O(N__3996),
            .I(ctrl_tap_fsm_state_2));
    LocalMux I__865 (
            .O(N__3987),
            .I(ctrl_tap_fsm_state_2));
    LocalMux I__864 (
            .O(N__3980),
            .I(ctrl_tap_fsm_state_2));
    LocalMux I__863 (
            .O(N__3973),
            .I(ctrl_tap_fsm_state_2));
    CascadeMux I__862 (
            .O(N__3956),
            .I(N__3946));
    CascadeMux I__861 (
            .O(N__3955),
            .I(N__3940));
    InMux I__860 (
            .O(N__3954),
            .I(N__3934));
    InMux I__859 (
            .O(N__3953),
            .I(N__3934));
    InMux I__858 (
            .O(N__3952),
            .I(N__3931));
    InMux I__857 (
            .O(N__3951),
            .I(N__3926));
    InMux I__856 (
            .O(N__3950),
            .I(N__3926));
    CascadeMux I__855 (
            .O(N__3949),
            .I(N__3923));
    InMux I__854 (
            .O(N__3946),
            .I(N__3920));
    InMux I__853 (
            .O(N__3945),
            .I(N__3913));
    InMux I__852 (
            .O(N__3944),
            .I(N__3913));
    InMux I__851 (
            .O(N__3943),
            .I(N__3913));
    InMux I__850 (
            .O(N__3940),
            .I(N__3907));
    InMux I__849 (
            .O(N__3939),
            .I(N__3907));
    LocalMux I__848 (
            .O(N__3934),
            .I(N__3900));
    LocalMux I__847 (
            .O(N__3931),
            .I(N__3900));
    LocalMux I__846 (
            .O(N__3926),
            .I(N__3900));
    InMux I__845 (
            .O(N__3923),
            .I(N__3897));
    LocalMux I__844 (
            .O(N__3920),
            .I(N__3892));
    LocalMux I__843 (
            .O(N__3913),
            .I(N__3892));
    InMux I__842 (
            .O(N__3912),
            .I(N__3889));
    LocalMux I__841 (
            .O(N__3907),
            .I(N__3886));
    Span4Mux_h I__840 (
            .O(N__3900),
            .I(N__3883));
    LocalMux I__839 (
            .O(N__3897),
            .I(N__3880));
    Span4Mux_h I__838 (
            .O(N__3892),
            .I(N__3877));
    LocalMux I__837 (
            .O(N__3889),
            .I(N__3874));
    Span12Mux_s8_h I__836 (
            .O(N__3886),
            .I(N__3871));
    Span4Mux_v I__835 (
            .O(N__3883),
            .I(N__3868));
    Span4Mux_h I__834 (
            .O(N__3880),
            .I(N__3865));
    Span4Mux_v I__833 (
            .O(N__3877),
            .I(N__3860));
    Span4Mux_v I__832 (
            .O(N__3874),
            .I(N__3860));
    Odrv12 I__831 (
            .O(N__3871),
            .I(ctrl_tap_fsm_stateNext_3__N_10_c_3));
    Odrv4 I__830 (
            .O(N__3868),
            .I(ctrl_tap_fsm_stateNext_3__N_10_c_3));
    Odrv4 I__829 (
            .O(N__3865),
            .I(ctrl_tap_fsm_stateNext_3__N_10_c_3));
    Odrv4 I__828 (
            .O(N__3860),
            .I(ctrl_tap_fsm_stateNext_3__N_10_c_3));
    CascadeMux I__827 (
            .O(N__3851),
            .I(N__3844));
    InMux I__826 (
            .O(N__3850),
            .I(N__3829));
    InMux I__825 (
            .O(N__3849),
            .I(N__3829));
    InMux I__824 (
            .O(N__3848),
            .I(N__3829));
    InMux I__823 (
            .O(N__3847),
            .I(N__3826));
    InMux I__822 (
            .O(N__3844),
            .I(N__3823));
    InMux I__821 (
            .O(N__3843),
            .I(N__3807));
    InMux I__820 (
            .O(N__3842),
            .I(N__3807));
    InMux I__819 (
            .O(N__3841),
            .I(N__3807));
    InMux I__818 (
            .O(N__3840),
            .I(N__3804));
    InMux I__817 (
            .O(N__3839),
            .I(N__3799));
    InMux I__816 (
            .O(N__3838),
            .I(N__3799));
    InMux I__815 (
            .O(N__3837),
            .I(N__3794));
    InMux I__814 (
            .O(N__3836),
            .I(N__3794));
    LocalMux I__813 (
            .O(N__3829),
            .I(N__3791));
    LocalMux I__812 (
            .O(N__3826),
            .I(N__3786));
    LocalMux I__811 (
            .O(N__3823),
            .I(N__3786));
    InMux I__810 (
            .O(N__3822),
            .I(N__3779));
    InMux I__809 (
            .O(N__3821),
            .I(N__3779));
    InMux I__808 (
            .O(N__3820),
            .I(N__3779));
    InMux I__807 (
            .O(N__3819),
            .I(N__3774));
    InMux I__806 (
            .O(N__3818),
            .I(N__3774));
    InMux I__805 (
            .O(N__3817),
            .I(N__3765));
    InMux I__804 (
            .O(N__3816),
            .I(N__3765));
    InMux I__803 (
            .O(N__3815),
            .I(N__3765));
    InMux I__802 (
            .O(N__3814),
            .I(N__3765));
    LocalMux I__801 (
            .O(N__3807),
            .I(ctrl_tap_fsm_state_1));
    LocalMux I__800 (
            .O(N__3804),
            .I(ctrl_tap_fsm_state_1));
    LocalMux I__799 (
            .O(N__3799),
            .I(ctrl_tap_fsm_state_1));
    LocalMux I__798 (
            .O(N__3794),
            .I(ctrl_tap_fsm_state_1));
    Odrv4 I__797 (
            .O(N__3791),
            .I(ctrl_tap_fsm_state_1));
    Odrv4 I__796 (
            .O(N__3786),
            .I(ctrl_tap_fsm_state_1));
    LocalMux I__795 (
            .O(N__3779),
            .I(ctrl_tap_fsm_state_1));
    LocalMux I__794 (
            .O(N__3774),
            .I(ctrl_tap_fsm_state_1));
    LocalMux I__793 (
            .O(N__3765),
            .I(ctrl_tap_fsm_state_1));
    InMux I__792 (
            .O(N__3746),
            .I(N__3743));
    LocalMux I__791 (
            .O(N__3743),
            .I(n2243));
    InMux I__790 (
            .O(N__3740),
            .I(N__3737));
    LocalMux I__789 (
            .O(N__3737),
            .I(n2186));
    InMux I__788 (
            .O(N__3734),
            .I(N__3727));
    CascadeMux I__787 (
            .O(N__3733),
            .I(N__3716));
    CascadeMux I__786 (
            .O(N__3732),
            .I(N__3712));
    InMux I__785 (
            .O(N__3731),
            .I(N__3708));
    CascadeMux I__784 (
            .O(N__3730),
            .I(N__3700));
    LocalMux I__783 (
            .O(N__3727),
            .I(N__3694));
    InMux I__782 (
            .O(N__3726),
            .I(N__3689));
    InMux I__781 (
            .O(N__3725),
            .I(N__3689));
    InMux I__780 (
            .O(N__3724),
            .I(N__3680));
    InMux I__779 (
            .O(N__3723),
            .I(N__3680));
    InMux I__778 (
            .O(N__3722),
            .I(N__3680));
    InMux I__777 (
            .O(N__3721),
            .I(N__3680));
    InMux I__776 (
            .O(N__3720),
            .I(N__3677));
    InMux I__775 (
            .O(N__3719),
            .I(N__3672));
    InMux I__774 (
            .O(N__3716),
            .I(N__3672));
    InMux I__773 (
            .O(N__3715),
            .I(N__3669));
    InMux I__772 (
            .O(N__3712),
            .I(N__3664));
    InMux I__771 (
            .O(N__3711),
            .I(N__3664));
    LocalMux I__770 (
            .O(N__3708),
            .I(N__3661));
    InMux I__769 (
            .O(N__3707),
            .I(N__3656));
    InMux I__768 (
            .O(N__3706),
            .I(N__3656));
    InMux I__767 (
            .O(N__3705),
            .I(N__3649));
    InMux I__766 (
            .O(N__3704),
            .I(N__3649));
    InMux I__765 (
            .O(N__3703),
            .I(N__3649));
    InMux I__764 (
            .O(N__3700),
            .I(N__3644));
    InMux I__763 (
            .O(N__3699),
            .I(N__3644));
    InMux I__762 (
            .O(N__3698),
            .I(N__3639));
    InMux I__761 (
            .O(N__3697),
            .I(N__3639));
    Odrv4 I__760 (
            .O(N__3694),
            .I(ctrl_tap_fsm_state_0));
    LocalMux I__759 (
            .O(N__3689),
            .I(ctrl_tap_fsm_state_0));
    LocalMux I__758 (
            .O(N__3680),
            .I(ctrl_tap_fsm_state_0));
    LocalMux I__757 (
            .O(N__3677),
            .I(ctrl_tap_fsm_state_0));
    LocalMux I__756 (
            .O(N__3672),
            .I(ctrl_tap_fsm_state_0));
    LocalMux I__755 (
            .O(N__3669),
            .I(ctrl_tap_fsm_state_0));
    LocalMux I__754 (
            .O(N__3664),
            .I(ctrl_tap_fsm_state_0));
    Odrv4 I__753 (
            .O(N__3661),
            .I(ctrl_tap_fsm_state_0));
    LocalMux I__752 (
            .O(N__3656),
            .I(ctrl_tap_fsm_state_0));
    LocalMux I__751 (
            .O(N__3649),
            .I(ctrl_tap_fsm_state_0));
    LocalMux I__750 (
            .O(N__3644),
            .I(ctrl_tap_fsm_state_0));
    LocalMux I__749 (
            .O(N__3639),
            .I(ctrl_tap_fsm_state_0));
    CascadeMux I__748 (
            .O(N__3614),
            .I(n17_cascade_));
    CascadeMux I__747 (
            .O(N__3611),
            .I(n1687_cascade_));
    InMux I__746 (
            .O(N__3608),
            .I(N__3605));
    LocalMux I__745 (
            .O(N__3605),
            .I(n2234));
    InMux I__744 (
            .O(N__3602),
            .I(N__3599));
    LocalMux I__743 (
            .O(N__3599),
            .I(n8));
    InMux I__742 (
            .O(N__3596),
            .I(N__3593));
    LocalMux I__741 (
            .O(N__3593),
            .I(n2198));
    InMux I__740 (
            .O(N__3590),
            .I(N__3586));
    InMux I__739 (
            .O(N__3589),
            .I(N__3583));
    LocalMux I__738 (
            .O(N__3586),
            .I(N__3580));
    LocalMux I__737 (
            .O(N__3583),
            .I(ctrl_tap_instructionShift_0));
    Odrv12 I__736 (
            .O(N__3580),
            .I(ctrl_tap_instructionShift_0));
    InMux I__735 (
            .O(N__3575),
            .I(N__3572));
    LocalMux I__734 (
            .O(N__3572),
            .I(ctrl_tap_bypass));
    CascadeMux I__733 (
            .O(N__3569),
            .I(n2198_cascade_));
    InMux I__732 (
            .O(N__3566),
            .I(N__3563));
    LocalMux I__731 (
            .O(N__3563),
            .I(n4));
    InMux I__730 (
            .O(N__3560),
            .I(N__3557));
    LocalMux I__729 (
            .O(N__3557),
            .I(ctrl_tap_tdoUnbufferd_N_213));
    CascadeMux I__728 (
            .O(N__3554),
            .I(N__3551));
    InMux I__727 (
            .O(N__3551),
            .I(N__3547));
    InMux I__726 (
            .O(N__3550),
            .I(N__3544));
    LocalMux I__725 (
            .O(N__3547),
            .I(ctrl_idcodeArea_shifter_27));
    LocalMux I__724 (
            .O(N__3544),
            .I(ctrl_idcodeArea_shifter_27));
    CascadeMux I__723 (
            .O(N__3539),
            .I(N__3535));
    CascadeMux I__722 (
            .O(N__3538),
            .I(N__3532));
    InMux I__721 (
            .O(N__3535),
            .I(N__3527));
    InMux I__720 (
            .O(N__3532),
            .I(N__3527));
    LocalMux I__719 (
            .O(N__3527),
            .I(ctrl_idcodeArea_shifter_26));
    InMux I__718 (
            .O(N__3524),
            .I(N__3519));
    InMux I__717 (
            .O(N__3523),
            .I(N__3516));
    InMux I__716 (
            .O(N__3522),
            .I(N__3513));
    LocalMux I__715 (
            .O(N__3519),
            .I(N__3509));
    LocalMux I__714 (
            .O(N__3516),
            .I(N__3506));
    LocalMux I__713 (
            .O(N__3513),
            .I(N__3503));
    InMux I__712 (
            .O(N__3512),
            .I(N__3500));
    Span4Mux_v I__711 (
            .O(N__3509),
            .I(N__3495));
    Span4Mux_h I__710 (
            .O(N__3506),
            .I(N__3495));
    Span4Mux_v I__709 (
            .O(N__3503),
            .I(N__3490));
    LocalMux I__708 (
            .O(N__3500),
            .I(N__3490));
    Odrv4 I__707 (
            .O(N__3495),
            .I(io_jtag_tdi_c));
    Odrv4 I__706 (
            .O(N__3490),
            .I(io_jtag_tdi_c));
    CascadeMux I__705 (
            .O(N__3485),
            .I(N__3481));
    InMux I__704 (
            .O(N__3484),
            .I(N__3478));
    InMux I__703 (
            .O(N__3481),
            .I(N__3475));
    LocalMux I__702 (
            .O(N__3478),
            .I(ctrl_idcodeArea_shifter_23));
    LocalMux I__701 (
            .O(N__3475),
            .I(ctrl_idcodeArea_shifter_23));
    CascadeMux I__700 (
            .O(N__3470),
            .I(N__3466));
    InMux I__699 (
            .O(N__3469),
            .I(N__3463));
    InMux I__698 (
            .O(N__3466),
            .I(N__3460));
    LocalMux I__697 (
            .O(N__3463),
            .I(ctrl_idcodeArea_shifter_22));
    LocalMux I__696 (
            .O(N__3460),
            .I(ctrl_idcodeArea_shifter_22));
    InMux I__695 (
            .O(N__3455),
            .I(N__3449));
    InMux I__694 (
            .O(N__3454),
            .I(N__3449));
    LocalMux I__693 (
            .O(N__3449),
            .I(ctrl_idcodeArea_shifter_21));
    CascadeMux I__692 (
            .O(N__3446),
            .I(N__3442));
    InMux I__691 (
            .O(N__3445),
            .I(N__3439));
    InMux I__690 (
            .O(N__3442),
            .I(N__3436));
    LocalMux I__689 (
            .O(N__3439),
            .I(ctrl_idcodeArea_shifter_18));
    LocalMux I__688 (
            .O(N__3436),
            .I(ctrl_idcodeArea_shifter_18));
    CascadeMux I__687 (
            .O(N__3431),
            .I(N__3397));
    InMux I__686 (
            .O(N__3430),
            .I(N__3388));
    InMux I__685 (
            .O(N__3429),
            .I(N__3388));
    InMux I__684 (
            .O(N__3428),
            .I(N__3388));
    InMux I__683 (
            .O(N__3427),
            .I(N__3388));
    InMux I__682 (
            .O(N__3426),
            .I(N__3371));
    InMux I__681 (
            .O(N__3425),
            .I(N__3371));
    InMux I__680 (
            .O(N__3424),
            .I(N__3371));
    InMux I__679 (
            .O(N__3423),
            .I(N__3371));
    InMux I__678 (
            .O(N__3422),
            .I(N__3371));
    InMux I__677 (
            .O(N__3421),
            .I(N__3371));
    InMux I__676 (
            .O(N__3420),
            .I(N__3371));
    InMux I__675 (
            .O(N__3419),
            .I(N__3371));
    InMux I__674 (
            .O(N__3418),
            .I(N__3360));
    InMux I__673 (
            .O(N__3417),
            .I(N__3360));
    InMux I__672 (
            .O(N__3416),
            .I(N__3360));
    InMux I__671 (
            .O(N__3415),
            .I(N__3360));
    InMux I__670 (
            .O(N__3414),
            .I(N__3360));
    InMux I__669 (
            .O(N__3413),
            .I(N__3349));
    InMux I__668 (
            .O(N__3412),
            .I(N__3349));
    InMux I__667 (
            .O(N__3411),
            .I(N__3349));
    InMux I__666 (
            .O(N__3410),
            .I(N__3349));
    InMux I__665 (
            .O(N__3409),
            .I(N__3349));
    InMux I__664 (
            .O(N__3408),
            .I(N__3332));
    InMux I__663 (
            .O(N__3407),
            .I(N__3332));
    InMux I__662 (
            .O(N__3406),
            .I(N__3332));
    InMux I__661 (
            .O(N__3405),
            .I(N__3332));
    InMux I__660 (
            .O(N__3404),
            .I(N__3332));
    InMux I__659 (
            .O(N__3403),
            .I(N__3332));
    InMux I__658 (
            .O(N__3402),
            .I(N__3332));
    InMux I__657 (
            .O(N__3401),
            .I(N__3332));
    InMux I__656 (
            .O(N__3400),
            .I(N__3327));
    InMux I__655 (
            .O(N__3397),
            .I(N__3327));
    LocalMux I__654 (
            .O(N__3388),
            .I(n15));
    LocalMux I__653 (
            .O(N__3371),
            .I(n15));
    LocalMux I__652 (
            .O(N__3360),
            .I(n15));
    LocalMux I__651 (
            .O(N__3349),
            .I(n15));
    LocalMux I__650 (
            .O(N__3332),
            .I(n15));
    LocalMux I__649 (
            .O(N__3327),
            .I(n15));
    CascadeMux I__648 (
            .O(N__3314),
            .I(N__3310));
    CascadeMux I__647 (
            .O(N__3313),
            .I(N__3307));
    InMux I__646 (
            .O(N__3310),
            .I(N__3302));
    InMux I__645 (
            .O(N__3307),
            .I(N__3302));
    LocalMux I__644 (
            .O(N__3302),
            .I(ctrl_idcodeArea_shifter_20));
    CascadeMux I__643 (
            .O(N__3299),
            .I(N__3287));
    CascadeMux I__642 (
            .O(N__3298),
            .I(N__3282));
    CascadeMux I__641 (
            .O(N__3297),
            .I(N__3279));
    CascadeMux I__640 (
            .O(N__3296),
            .I(N__3275));
    CascadeMux I__639 (
            .O(N__3295),
            .I(N__3272));
    CascadeMux I__638 (
            .O(N__3294),
            .I(N__3267));
    CascadeMux I__637 (
            .O(N__3293),
            .I(N__3263));
    CascadeMux I__636 (
            .O(N__3292),
            .I(N__3260));
    InMux I__635 (
            .O(N__3291),
            .I(N__3250));
    InMux I__634 (
            .O(N__3290),
            .I(N__3250));
    InMux I__633 (
            .O(N__3287),
            .I(N__3250));
    InMux I__632 (
            .O(N__3286),
            .I(N__3250));
    InMux I__631 (
            .O(N__3285),
            .I(N__3220));
    InMux I__630 (
            .O(N__3282),
            .I(N__3220));
    InMux I__629 (
            .O(N__3279),
            .I(N__3220));
    InMux I__628 (
            .O(N__3278),
            .I(N__3220));
    InMux I__627 (
            .O(N__3275),
            .I(N__3220));
    InMux I__626 (
            .O(N__3272),
            .I(N__3220));
    InMux I__625 (
            .O(N__3271),
            .I(N__3220));
    InMux I__624 (
            .O(N__3270),
            .I(N__3220));
    InMux I__623 (
            .O(N__3267),
            .I(N__3209));
    InMux I__622 (
            .O(N__3266),
            .I(N__3209));
    InMux I__621 (
            .O(N__3263),
            .I(N__3209));
    InMux I__620 (
            .O(N__3260),
            .I(N__3209));
    InMux I__619 (
            .O(N__3259),
            .I(N__3209));
    LocalMux I__618 (
            .O(N__3250),
            .I(N__3200));
    InMux I__617 (
            .O(N__3249),
            .I(N__3193));
    InMux I__616 (
            .O(N__3248),
            .I(N__3193));
    InMux I__615 (
            .O(N__3247),
            .I(N__3193));
    InMux I__614 (
            .O(N__3246),
            .I(N__3188));
    InMux I__613 (
            .O(N__3245),
            .I(N__3188));
    InMux I__612 (
            .O(N__3244),
            .I(N__3179));
    InMux I__611 (
            .O(N__3243),
            .I(N__3179));
    InMux I__610 (
            .O(N__3242),
            .I(N__3179));
    InMux I__609 (
            .O(N__3241),
            .I(N__3179));
    InMux I__608 (
            .O(N__3240),
            .I(N__3170));
    InMux I__607 (
            .O(N__3239),
            .I(N__3170));
    InMux I__606 (
            .O(N__3238),
            .I(N__3170));
    InMux I__605 (
            .O(N__3237),
            .I(N__3170));
    LocalMux I__604 (
            .O(N__3220),
            .I(N__3165));
    LocalMux I__603 (
            .O(N__3209),
            .I(N__3165));
    InMux I__602 (
            .O(N__3208),
            .I(N__3160));
    InMux I__601 (
            .O(N__3207),
            .I(N__3160));
    InMux I__600 (
            .O(N__3206),
            .I(N__3151));
    InMux I__599 (
            .O(N__3205),
            .I(N__3151));
    InMux I__598 (
            .O(N__3204),
            .I(N__3151));
    InMux I__597 (
            .O(N__3203),
            .I(N__3151));
    Odrv4 I__596 (
            .O(N__3200),
            .I(n1489));
    LocalMux I__595 (
            .O(N__3193),
            .I(n1489));
    LocalMux I__594 (
            .O(N__3188),
            .I(n1489));
    LocalMux I__593 (
            .O(N__3179),
            .I(n1489));
    LocalMux I__592 (
            .O(N__3170),
            .I(n1489));
    Odrv4 I__591 (
            .O(N__3165),
            .I(n1489));
    LocalMux I__590 (
            .O(N__3160),
            .I(n1489));
    LocalMux I__589 (
            .O(N__3151),
            .I(n1489));
    CascadeMux I__588 (
            .O(N__3134),
            .I(N__3130));
    InMux I__587 (
            .O(N__3133),
            .I(N__3125));
    InMux I__586 (
            .O(N__3130),
            .I(N__3125));
    LocalMux I__585 (
            .O(N__3125),
            .I(ctrl_idcodeArea_shifter_19));
    CascadeMux I__584 (
            .O(N__3122),
            .I(n2185_cascade_));
    InMux I__583 (
            .O(N__3119),
            .I(N__3099));
    InMux I__582 (
            .O(N__3118),
            .I(N__3099));
    InMux I__581 (
            .O(N__3117),
            .I(N__3099));
    InMux I__580 (
            .O(N__3116),
            .I(N__3099));
    InMux I__579 (
            .O(N__3115),
            .I(N__3079));
    InMux I__578 (
            .O(N__3114),
            .I(N__3079));
    InMux I__577 (
            .O(N__3113),
            .I(N__3079));
    InMux I__576 (
            .O(N__3112),
            .I(N__3079));
    InMux I__575 (
            .O(N__3111),
            .I(N__3070));
    InMux I__574 (
            .O(N__3110),
            .I(N__3070));
    InMux I__573 (
            .O(N__3109),
            .I(N__3070));
    InMux I__572 (
            .O(N__3108),
            .I(N__3070));
    LocalMux I__571 (
            .O(N__3099),
            .I(N__3067));
    InMux I__570 (
            .O(N__3098),
            .I(N__3058));
    InMux I__569 (
            .O(N__3097),
            .I(N__3058));
    InMux I__568 (
            .O(N__3096),
            .I(N__3058));
    InMux I__567 (
            .O(N__3095),
            .I(N__3058));
    InMux I__566 (
            .O(N__3094),
            .I(N__3051));
    InMux I__565 (
            .O(N__3093),
            .I(N__3051));
    InMux I__564 (
            .O(N__3092),
            .I(N__3051));
    InMux I__563 (
            .O(N__3091),
            .I(N__3042));
    InMux I__562 (
            .O(N__3090),
            .I(N__3042));
    InMux I__561 (
            .O(N__3089),
            .I(N__3042));
    InMux I__560 (
            .O(N__3088),
            .I(N__3042));
    LocalMux I__559 (
            .O(N__3079),
            .I(n1848));
    LocalMux I__558 (
            .O(N__3070),
            .I(n1848));
    Odrv4 I__557 (
            .O(N__3067),
            .I(n1848));
    LocalMux I__556 (
            .O(N__3058),
            .I(n1848));
    LocalMux I__555 (
            .O(N__3051),
            .I(n1848));
    LocalMux I__554 (
            .O(N__3042),
            .I(n1848));
    InMux I__553 (
            .O(N__3029),
            .I(N__3025));
    InMux I__552 (
            .O(N__3028),
            .I(N__3022));
    LocalMux I__551 (
            .O(N__3025),
            .I(myClockArea_timeout_counter_value_7));
    LocalMux I__550 (
            .O(N__3022),
            .I(myClockArea_timeout_counter_value_7));
    InMux I__549 (
            .O(N__3017),
            .I(N__3013));
    InMux I__548 (
            .O(N__3016),
            .I(N__3010));
    LocalMux I__547 (
            .O(N__3013),
            .I(myClockArea_timeout_counter_value_21));
    LocalMux I__546 (
            .O(N__3010),
            .I(myClockArea_timeout_counter_value_21));
    InMux I__545 (
            .O(N__3005),
            .I(N__3002));
    LocalMux I__544 (
            .O(N__3002),
            .I(n11));
    InMux I__543 (
            .O(N__2999),
            .I(N__2995));
    InMux I__542 (
            .O(N__2998),
            .I(N__2992));
    LocalMux I__541 (
            .O(N__2995),
            .I(myClockArea_timeout_counter_value_19));
    LocalMux I__540 (
            .O(N__2992),
            .I(myClockArea_timeout_counter_value_19));
    InMux I__539 (
            .O(N__2987),
            .I(N__2983));
    InMux I__538 (
            .O(N__2986),
            .I(N__2980));
    LocalMux I__537 (
            .O(N__2983),
            .I(myClockArea_timeout_counter_value_15));
    LocalMux I__536 (
            .O(N__2980),
            .I(myClockArea_timeout_counter_value_15));
    CascadeMux I__535 (
            .O(N__2975),
            .I(N__2971));
    InMux I__534 (
            .O(N__2974),
            .I(N__2968));
    InMux I__533 (
            .O(N__2971),
            .I(N__2965));
    LocalMux I__532 (
            .O(N__2968),
            .I(myClockArea_timeout_counter_value_20));
    LocalMux I__531 (
            .O(N__2965),
            .I(myClockArea_timeout_counter_value_20));
    InMux I__530 (
            .O(N__2960),
            .I(N__2956));
    InMux I__529 (
            .O(N__2959),
            .I(N__2953));
    LocalMux I__528 (
            .O(N__2956),
            .I(myClockArea_timeout_counter_value_11));
    LocalMux I__527 (
            .O(N__2953),
            .I(myClockArea_timeout_counter_value_11));
    InMux I__526 (
            .O(N__2948),
            .I(N__2945));
    LocalMux I__525 (
            .O(N__2945),
            .I(n2220));
    InMux I__524 (
            .O(N__2942),
            .I(N__2938));
    InMux I__523 (
            .O(N__2941),
            .I(N__2935));
    LocalMux I__522 (
            .O(N__2938),
            .I(myClockArea_timeout_counter_value_9));
    LocalMux I__521 (
            .O(N__2935),
            .I(myClockArea_timeout_counter_value_9));
    InMux I__520 (
            .O(N__2930),
            .I(N__2926));
    InMux I__519 (
            .O(N__2929),
            .I(N__2923));
    LocalMux I__518 (
            .O(N__2926),
            .I(myClockArea_timeout_counter_value_18));
    LocalMux I__517 (
            .O(N__2923),
            .I(myClockArea_timeout_counter_value_18));
    CascadeMux I__516 (
            .O(N__2918),
            .I(N__2914));
    InMux I__515 (
            .O(N__2917),
            .I(N__2911));
    InMux I__514 (
            .O(N__2914),
            .I(N__2908));
    LocalMux I__513 (
            .O(N__2911),
            .I(myClockArea_timeout_counter_value_12));
    LocalMux I__512 (
            .O(N__2908),
            .I(myClockArea_timeout_counter_value_12));
    InMux I__511 (
            .O(N__2903),
            .I(N__2899));
    InMux I__510 (
            .O(N__2902),
            .I(N__2896));
    LocalMux I__509 (
            .O(N__2899),
            .I(myClockArea_timeout_counter_value_14));
    LocalMux I__508 (
            .O(N__2896),
            .I(myClockArea_timeout_counter_value_14));
    InMux I__507 (
            .O(N__2891),
            .I(N__2888));
    LocalMux I__506 (
            .O(N__2888),
            .I(n13));
    InMux I__505 (
            .O(N__2885),
            .I(N__2880));
    InMux I__504 (
            .O(N__2884),
            .I(N__2877));
    InMux I__503 (
            .O(N__2883),
            .I(N__2874));
    LocalMux I__502 (
            .O(N__2880),
            .I(N__2871));
    LocalMux I__501 (
            .O(N__2877),
            .I(myClockArea_timeout_state));
    LocalMux I__500 (
            .O(N__2874),
            .I(myClockArea_timeout_state));
    Odrv4 I__499 (
            .O(N__2871),
            .I(myClockArea_timeout_state));
    IoInMux I__498 (
            .O(N__2864),
            .I(N__2861));
    LocalMux I__497 (
            .O(N__2861),
            .I(N__2857));
    InMux I__496 (
            .O(N__2860),
            .I(N__2854));
    Odrv12 I__495 (
            .O(N__2857),
            .I(io_leds_c_3));
    LocalMux I__494 (
            .O(N__2854),
            .I(io_leds_c_3));
    ClkMux I__493 (
            .O(N__2849),
            .I(N__2834));
    ClkMux I__492 (
            .O(N__2848),
            .I(N__2834));
    ClkMux I__491 (
            .O(N__2847),
            .I(N__2834));
    ClkMux I__490 (
            .O(N__2846),
            .I(N__2834));
    ClkMux I__489 (
            .O(N__2845),
            .I(N__2834));
    GlobalMux I__488 (
            .O(N__2834),
            .I(N__2831));
    gio2CtrlBuf I__487 (
            .O(N__2831),
            .I(global_clk_c));
    InMux I__486 (
            .O(N__2828),
            .I(N__2822));
    InMux I__485 (
            .O(N__2827),
            .I(N__2822));
    LocalMux I__484 (
            .O(N__2822),
            .I(ctrl_idcodeArea_shifter_25));
    CascadeMux I__483 (
            .O(N__2819),
            .I(N__2815));
    InMux I__482 (
            .O(N__2818),
            .I(N__2810));
    InMux I__481 (
            .O(N__2815),
            .I(N__2810));
    LocalMux I__480 (
            .O(N__2810),
            .I(ctrl_idcodeArea_shifter_24));
    IoInMux I__479 (
            .O(N__2807),
            .I(N__2804));
    LocalMux I__478 (
            .O(N__2804),
            .I(N__2801));
    IoSpan4Mux I__477 (
            .O(N__2801),
            .I(N__2797));
    CascadeMux I__476 (
            .O(N__2800),
            .I(N__2793));
    Span4Mux_s3_h I__475 (
            .O(N__2797),
            .I(N__2790));
    InMux I__474 (
            .O(N__2796),
            .I(N__2787));
    InMux I__473 (
            .O(N__2793),
            .I(N__2784));
    Odrv4 I__472 (
            .O(N__2790),
            .I(io_leds_c_7));
    LocalMux I__471 (
            .O(N__2787),
            .I(io_leds_c_7));
    LocalMux I__470 (
            .O(N__2784),
            .I(io_leds_c_7));
    InMux I__469 (
            .O(N__2777),
            .I(N__2773));
    InMux I__468 (
            .O(N__2776),
            .I(N__2770));
    LocalMux I__467 (
            .O(N__2773),
            .I(myClockArea_timeout_counter_value_3));
    LocalMux I__466 (
            .O(N__2770),
            .I(myClockArea_timeout_counter_value_3));
    InMux I__465 (
            .O(N__2765),
            .I(N__2761));
    InMux I__464 (
            .O(N__2764),
            .I(N__2758));
    LocalMux I__463 (
            .O(N__2761),
            .I(myClockArea_timeout_counter_value_1));
    LocalMux I__462 (
            .O(N__2758),
            .I(myClockArea_timeout_counter_value_1));
    CascadeMux I__461 (
            .O(N__2753),
            .I(N__2749));
    InMux I__460 (
            .O(N__2752),
            .I(N__2746));
    InMux I__459 (
            .O(N__2749),
            .I(N__2743));
    LocalMux I__458 (
            .O(N__2746),
            .I(myClockArea_timeout_counter_value_5));
    LocalMux I__457 (
            .O(N__2743),
            .I(myClockArea_timeout_counter_value_5));
    InMux I__456 (
            .O(N__2738),
            .I(N__2734));
    InMux I__455 (
            .O(N__2737),
            .I(N__2731));
    LocalMux I__454 (
            .O(N__2734),
            .I(myClockArea_timeout_counter_value_0));
    LocalMux I__453 (
            .O(N__2731),
            .I(myClockArea_timeout_counter_value_0));
    InMux I__452 (
            .O(N__2726),
            .I(N__2723));
    LocalMux I__451 (
            .O(N__2723),
            .I(n2309));
    InMux I__450 (
            .O(N__2720),
            .I(N__2716));
    InMux I__449 (
            .O(N__2719),
            .I(N__2713));
    LocalMux I__448 (
            .O(N__2716),
            .I(myClockArea_timeout_counter_value_4));
    LocalMux I__447 (
            .O(N__2713),
            .I(myClockArea_timeout_counter_value_4));
    InMux I__446 (
            .O(N__2708),
            .I(N__2704));
    InMux I__445 (
            .O(N__2707),
            .I(N__2701));
    LocalMux I__444 (
            .O(N__2704),
            .I(myClockArea_timeout_counter_value_6));
    LocalMux I__443 (
            .O(N__2701),
            .I(myClockArea_timeout_counter_value_6));
    CascadeMux I__442 (
            .O(N__2696),
            .I(N__2692));
    InMux I__441 (
            .O(N__2695),
            .I(N__2689));
    InMux I__440 (
            .O(N__2692),
            .I(N__2686));
    LocalMux I__439 (
            .O(N__2689),
            .I(myClockArea_timeout_counter_value_22));
    LocalMux I__438 (
            .O(N__2686),
            .I(myClockArea_timeout_counter_value_22));
    InMux I__437 (
            .O(N__2681),
            .I(N__2677));
    InMux I__436 (
            .O(N__2680),
            .I(N__2674));
    LocalMux I__435 (
            .O(N__2677),
            .I(myClockArea_timeout_counter_value_16));
    LocalMux I__434 (
            .O(N__2674),
            .I(myClockArea_timeout_counter_value_16));
    InMux I__433 (
            .O(N__2669),
            .I(N__2665));
    InMux I__432 (
            .O(N__2668),
            .I(N__2662));
    LocalMux I__431 (
            .O(N__2665),
            .I(myClockArea_timeout_counter_value_17));
    LocalMux I__430 (
            .O(N__2662),
            .I(myClockArea_timeout_counter_value_17));
    InMux I__429 (
            .O(N__2657),
            .I(N__2653));
    InMux I__428 (
            .O(N__2656),
            .I(N__2650));
    LocalMux I__427 (
            .O(N__2653),
            .I(myClockArea_timeout_counter_value_8));
    LocalMux I__426 (
            .O(N__2650),
            .I(myClockArea_timeout_counter_value_8));
    CascadeMux I__425 (
            .O(N__2645),
            .I(N__2641));
    InMux I__424 (
            .O(N__2644),
            .I(N__2638));
    InMux I__423 (
            .O(N__2641),
            .I(N__2635));
    LocalMux I__422 (
            .O(N__2638),
            .I(myClockArea_timeout_counter_value_10));
    LocalMux I__421 (
            .O(N__2635),
            .I(myClockArea_timeout_counter_value_10));
    InMux I__420 (
            .O(N__2630),
            .I(N__2626));
    InMux I__419 (
            .O(N__2629),
            .I(N__2623));
    LocalMux I__418 (
            .O(N__2626),
            .I(myClockArea_timeout_counter_value_2));
    LocalMux I__417 (
            .O(N__2623),
            .I(myClockArea_timeout_counter_value_2));
    InMux I__416 (
            .O(N__2618),
            .I(N__2615));
    LocalMux I__415 (
            .O(N__2615),
            .I(n2216));
    CascadeMux I__414 (
            .O(N__2612),
            .I(n2218_cascade_));
    InMux I__413 (
            .O(N__2609),
            .I(N__2606));
    LocalMux I__412 (
            .O(N__2606),
            .I(n2222));
    InMux I__411 (
            .O(N__2603),
            .I(N__2599));
    InMux I__410 (
            .O(N__2602),
            .I(N__2596));
    LocalMux I__409 (
            .O(N__2599),
            .I(myClockArea_timeout_counter_value_13));
    LocalMux I__408 (
            .O(N__2596),
            .I(myClockArea_timeout_counter_value_13));
    CascadeMux I__407 (
            .O(N__2591),
            .I(n2228_cascade_));
    InMux I__406 (
            .O(N__2588),
            .I(N__2585));
    LocalMux I__405 (
            .O(N__2585),
            .I(N__2582));
    Odrv4 I__404 (
            .O(N__2582),
            .I(n2185));
    CascadeMux I__403 (
            .O(N__2579),
            .I(n2282_cascade_));
    CascadeMux I__402 (
            .O(N__2576),
            .I(n2326_cascade_));
    InMux I__401 (
            .O(N__2573),
            .I(N__2570));
    LocalMux I__400 (
            .O(N__2570),
            .I(n2306));
    CascadeMux I__399 (
            .O(N__2567),
            .I(N__2563));
    CEMux I__398 (
            .O(N__2566),
            .I(N__2560));
    InMux I__397 (
            .O(N__2563),
            .I(N__2557));
    LocalMux I__396 (
            .O(N__2560),
            .I(n1022));
    LocalMux I__395 (
            .O(N__2557),
            .I(n1022));
    CascadeMux I__394 (
            .O(N__2552),
            .I(n2231_cascade_));
    InMux I__393 (
            .O(N__2549),
            .I(N__2546));
    LocalMux I__392 (
            .O(N__2546),
            .I(n2273));
    CascadeMux I__391 (
            .O(N__2543),
            .I(n2263_cascade_));
    InMux I__390 (
            .O(N__2540),
            .I(N__2537));
    LocalMux I__389 (
            .O(N__2537),
            .I(n2323));
    InMux I__388 (
            .O(N__2534),
            .I(N__2531));
    LocalMux I__387 (
            .O(N__2531),
            .I(n2272));
    CascadeMux I__386 (
            .O(N__2528),
            .I(n1489_cascade_));
    CascadeMux I__385 (
            .O(N__2525),
            .I(n1269_cascade_));
    InMux I__384 (
            .O(N__2522),
            .I(N__2515));
    InMux I__383 (
            .O(N__2521),
            .I(N__2512));
    InMux I__382 (
            .O(N__2520),
            .I(N__2509));
    InMux I__381 (
            .O(N__2519),
            .I(N__2504));
    InMux I__380 (
            .O(N__2518),
            .I(N__2504));
    LocalMux I__379 (
            .O(N__2515),
            .I(ctrl_tap_instruction_0));
    LocalMux I__378 (
            .O(N__2512),
            .I(ctrl_tap_instruction_0));
    LocalMux I__377 (
            .O(N__2509),
            .I(ctrl_tap_instruction_0));
    LocalMux I__376 (
            .O(N__2504),
            .I(ctrl_tap_instruction_0));
    CascadeMux I__375 (
            .O(N__2495),
            .I(N__2492));
    InMux I__374 (
            .O(N__2492),
            .I(N__2488));
    InMux I__373 (
            .O(N__2491),
            .I(N__2485));
    LocalMux I__372 (
            .O(N__2488),
            .I(ctrl_tap_instructionShift_3));
    LocalMux I__371 (
            .O(N__2485),
            .I(ctrl_tap_instructionShift_3));
    InMux I__370 (
            .O(N__2480),
            .I(N__2476));
    CascadeMux I__369 (
            .O(N__2479),
            .I(N__2471));
    LocalMux I__368 (
            .O(N__2476),
            .I(N__2467));
    InMux I__367 (
            .O(N__2475),
            .I(N__2464));
    InMux I__366 (
            .O(N__2474),
            .I(N__2461));
    InMux I__365 (
            .O(N__2471),
            .I(N__2456));
    InMux I__364 (
            .O(N__2470),
            .I(N__2456));
    Odrv4 I__363 (
            .O(N__2467),
            .I(ctrl_tap_instruction_3));
    LocalMux I__362 (
            .O(N__2464),
            .I(ctrl_tap_instruction_3));
    LocalMux I__361 (
            .O(N__2461),
            .I(ctrl_tap_instruction_3));
    LocalMux I__360 (
            .O(N__2456),
            .I(ctrl_tap_instruction_3));
    CascadeMux I__359 (
            .O(N__2447),
            .I(N__2444));
    InMux I__358 (
            .O(N__2444),
            .I(N__2440));
    InMux I__357 (
            .O(N__2443),
            .I(N__2437));
    LocalMux I__356 (
            .O(N__2440),
            .I(ctrl_tap_instructionShift_2));
    LocalMux I__355 (
            .O(N__2437),
            .I(ctrl_tap_instructionShift_2));
    InMux I__354 (
            .O(N__2432),
            .I(N__2425));
    InMux I__353 (
            .O(N__2431),
            .I(N__2422));
    InMux I__352 (
            .O(N__2430),
            .I(N__2419));
    InMux I__351 (
            .O(N__2429),
            .I(N__2414));
    InMux I__350 (
            .O(N__2428),
            .I(N__2414));
    LocalMux I__349 (
            .O(N__2425),
            .I(ctrl_tap_instruction_2));
    LocalMux I__348 (
            .O(N__2422),
            .I(ctrl_tap_instruction_2));
    LocalMux I__347 (
            .O(N__2419),
            .I(ctrl_tap_instruction_2));
    LocalMux I__346 (
            .O(N__2414),
            .I(ctrl_tap_instruction_2));
    InMux I__345 (
            .O(N__2405),
            .I(N__2396));
    InMux I__344 (
            .O(N__2404),
            .I(N__2396));
    InMux I__343 (
            .O(N__2403),
            .I(N__2396));
    LocalMux I__342 (
            .O(N__2396),
            .I(n1269));
    CascadeMux I__341 (
            .O(N__2393),
            .I(N__2390));
    InMux I__340 (
            .O(N__2390),
            .I(N__2386));
    InMux I__339 (
            .O(N__2389),
            .I(N__2383));
    LocalMux I__338 (
            .O(N__2386),
            .I(ctrl_tap_instructionShift_1));
    LocalMux I__337 (
            .O(N__2383),
            .I(ctrl_tap_instructionShift_1));
    CascadeMux I__336 (
            .O(N__2378),
            .I(N__2373));
    InMux I__335 (
            .O(N__2377),
            .I(N__2368));
    InMux I__334 (
            .O(N__2376),
            .I(N__2365));
    InMux I__333 (
            .O(N__2373),
            .I(N__2362));
    InMux I__332 (
            .O(N__2372),
            .I(N__2359));
    InMux I__331 (
            .O(N__2371),
            .I(N__2356));
    LocalMux I__330 (
            .O(N__2368),
            .I(ctrl_tap_instruction_1));
    LocalMux I__329 (
            .O(N__2365),
            .I(ctrl_tap_instruction_1));
    LocalMux I__328 (
            .O(N__2362),
            .I(ctrl_tap_instruction_1));
    LocalMux I__327 (
            .O(N__2359),
            .I(ctrl_tap_instruction_1));
    LocalMux I__326 (
            .O(N__2356),
            .I(ctrl_tap_instruction_1));
    InMux I__325 (
            .O(N__2345),
            .I(N__2342));
    LocalMux I__324 (
            .O(N__2342),
            .I(n2248));
    CascadeMux I__323 (
            .O(N__2339),
            .I(n118_cascade_));
    CascadeMux I__322 (
            .O(N__2336),
            .I(N__2333));
    InMux I__321 (
            .O(N__2333),
            .I(N__2329));
    InMux I__320 (
            .O(N__2332),
            .I(N__2326));
    LocalMux I__319 (
            .O(N__2329),
            .I(N__2323));
    LocalMux I__318 (
            .O(N__2326),
            .I(ctrl_idcodeArea_shifter_17));
    Odrv12 I__317 (
            .O(N__2323),
            .I(ctrl_idcodeArea_shifter_17));
    InMux I__316 (
            .O(N__2318),
            .I(N__2314));
    InMux I__315 (
            .O(N__2317),
            .I(N__2311));
    LocalMux I__314 (
            .O(N__2314),
            .I(ctrl_idcodeArea_shifter_1));
    LocalMux I__313 (
            .O(N__2311),
            .I(ctrl_idcodeArea_shifter_1));
    CascadeMux I__312 (
            .O(N__2306),
            .I(n6_cascade_));
    InMux I__311 (
            .O(N__2303),
            .I(N__2297));
    InMux I__310 (
            .O(N__2302),
            .I(N__2297));
    LocalMux I__309 (
            .O(N__2297),
            .I(ctrl_idcodeArea_shifter_0));
    InMux I__308 (
            .O(N__2294),
            .I(N__2291));
    LocalMux I__307 (
            .O(N__2291),
            .I(n2085));
    CascadeMux I__306 (
            .O(N__2288),
            .I(n15_cascade_));
    CascadeMux I__305 (
            .O(N__2285),
            .I(N__2281));
    InMux I__304 (
            .O(N__2284),
            .I(N__2278));
    InMux I__303 (
            .O(N__2281),
            .I(N__2275));
    LocalMux I__302 (
            .O(N__2278),
            .I(N__2272));
    LocalMux I__301 (
            .O(N__2275),
            .I(n7_adj_1));
    Odrv4 I__300 (
            .O(N__2272),
            .I(n7_adj_1));
    InMux I__299 (
            .O(N__2267),
            .I(N__2264));
    LocalMux I__298 (
            .O(N__2264),
            .I(N__2260));
    InMux I__297 (
            .O(N__2263),
            .I(N__2257));
    Span4Mux_h I__296 (
            .O(N__2260),
            .I(N__2254));
    LocalMux I__295 (
            .O(N__2257),
            .I(ctrl_ledsArea_shifter_0));
    Odrv4 I__294 (
            .O(N__2254),
            .I(ctrl_ledsArea_shifter_0));
    CascadeMux I__293 (
            .O(N__2249),
            .I(ctrl_tap_tdoUnbufferd_N_211_cascade_));
    IoInMux I__292 (
            .O(N__2246),
            .I(N__2243));
    LocalMux I__291 (
            .O(N__2243),
            .I(N__2240));
    Odrv12 I__290 (
            .O(N__2240),
            .I(ctrl_tap_tdoUnbufferd));
    InMux I__289 (
            .O(N__2237),
            .I(n2078));
    InMux I__288 (
            .O(N__2234),
            .I(n2079));
    InMux I__287 (
            .O(N__2231),
            .I(n2080));
    SRMux I__286 (
            .O(N__2228),
            .I(N__2224));
    SRMux I__285 (
            .O(N__2227),
            .I(N__2220));
    LocalMux I__284 (
            .O(N__2224),
            .I(N__2217));
    SRMux I__283 (
            .O(N__2223),
            .I(N__2214));
    LocalMux I__282 (
            .O(N__2220),
            .I(N__2210));
    Span4Mux_v I__281 (
            .O(N__2217),
            .I(N__2205));
    LocalMux I__280 (
            .O(N__2214),
            .I(N__2205));
    SRMux I__279 (
            .O(N__2213),
            .I(N__2202));
    Span4Mux_v I__278 (
            .O(N__2210),
            .I(N__2195));
    Span4Mux_h I__277 (
            .O(N__2205),
            .I(N__2195));
    LocalMux I__276 (
            .O(N__2202),
            .I(N__2195));
    Span4Mux_v I__275 (
            .O(N__2195),
            .I(N__2192));
    IoSpan4Mux I__274 (
            .O(N__2192),
            .I(N__2189));
    Odrv4 I__273 (
            .O(N__2189),
            .I(global_reset_c));
    InMux I__272 (
            .O(N__2186),
            .I(N__2180));
    InMux I__271 (
            .O(N__2185),
            .I(N__2180));
    LocalMux I__270 (
            .O(N__2180),
            .I(ctrl_idcodeArea_shifter_31));
    InMux I__269 (
            .O(N__2177),
            .I(N__2171));
    InMux I__268 (
            .O(N__2176),
            .I(N__2171));
    LocalMux I__267 (
            .O(N__2171),
            .I(ctrl_idcodeArea_shifter_28));
    CascadeMux I__266 (
            .O(N__2168),
            .I(N__2165));
    InMux I__265 (
            .O(N__2165),
            .I(N__2159));
    InMux I__264 (
            .O(N__2164),
            .I(N__2159));
    LocalMux I__263 (
            .O(N__2159),
            .I(ctrl_idcodeArea_shifter_30));
    InMux I__262 (
            .O(N__2156),
            .I(N__2150));
    InMux I__261 (
            .O(N__2155),
            .I(N__2150));
    LocalMux I__260 (
            .O(N__2150),
            .I(ctrl_idcodeArea_shifter_29));
    InMux I__259 (
            .O(N__2147),
            .I(n2069));
    InMux I__258 (
            .O(N__2144),
            .I(n2070));
    InMux I__257 (
            .O(N__2141),
            .I(n2071));
    InMux I__256 (
            .O(N__2138),
            .I(n2072));
    InMux I__255 (
            .O(N__2135),
            .I(n2073));
    InMux I__254 (
            .O(N__2132),
            .I(bfn_4_9_0_));
    InMux I__253 (
            .O(N__2129),
            .I(n2075));
    InMux I__252 (
            .O(N__2126),
            .I(n2076));
    InMux I__251 (
            .O(N__2123),
            .I(n2077));
    InMux I__250 (
            .O(N__2120),
            .I(n2060));
    InMux I__249 (
            .O(N__2117),
            .I(n2061));
    InMux I__248 (
            .O(N__2114),
            .I(n2062));
    InMux I__247 (
            .O(N__2111),
            .I(n2063));
    InMux I__246 (
            .O(N__2108),
            .I(n2064));
    InMux I__245 (
            .O(N__2105),
            .I(n2065));
    InMux I__244 (
            .O(N__2102),
            .I(bfn_4_8_0_));
    InMux I__243 (
            .O(N__2099),
            .I(n2067));
    InMux I__242 (
            .O(N__2096),
            .I(n2068));
    InMux I__241 (
            .O(N__2093),
            .I(N__2090));
    LocalMux I__240 (
            .O(N__2090),
            .I(N__2087));
    Odrv4 I__239 (
            .O(N__2087),
            .I(n7));
    CascadeMux I__238 (
            .O(N__2084),
            .I(n7_cascade_));
    InMux I__237 (
            .O(N__2081),
            .I(N__2078));
    LocalMux I__236 (
            .O(N__2078),
            .I(n2206));
    CascadeMux I__235 (
            .O(N__2075),
            .I(n7_adj_1_cascade_));
    InMux I__234 (
            .O(N__2072),
            .I(bfn_4_7_0_));
    InMux I__233 (
            .O(N__2069),
            .I(n2059));
    InMux I__232 (
            .O(N__2066),
            .I(N__2060));
    InMux I__231 (
            .O(N__2065),
            .I(N__2060));
    LocalMux I__230 (
            .O(N__2060),
            .I(ctrl_idcodeArea_shifter_16));
    CascadeMux I__229 (
            .O(N__2057),
            .I(N__2053));
    CascadeMux I__228 (
            .O(N__2056),
            .I(N__2050));
    InMux I__227 (
            .O(N__2053),
            .I(N__2045));
    InMux I__226 (
            .O(N__2050),
            .I(N__2045));
    LocalMux I__225 (
            .O(N__2045),
            .I(ctrl_idcodeArea_shifter_15));
    CascadeMux I__224 (
            .O(N__2042),
            .I(N__2038));
    InMux I__223 (
            .O(N__2041),
            .I(N__2033));
    InMux I__222 (
            .O(N__2038),
            .I(N__2033));
    LocalMux I__221 (
            .O(N__2033),
            .I(ctrl_idcodeArea_shifter_14));
    CascadeMux I__220 (
            .O(N__2030),
            .I(N__2026));
    InMux I__219 (
            .O(N__2029),
            .I(N__2021));
    InMux I__218 (
            .O(N__2026),
            .I(N__2021));
    LocalMux I__217 (
            .O(N__2021),
            .I(ctrl_idcodeArea_shifter_13));
    CascadeMux I__216 (
            .O(N__2018),
            .I(N__2014));
    InMux I__215 (
            .O(N__2017),
            .I(N__2009));
    InMux I__214 (
            .O(N__2014),
            .I(N__2009));
    LocalMux I__213 (
            .O(N__2009),
            .I(ctrl_idcodeArea_shifter_12));
    CascadeMux I__212 (
            .O(N__2006),
            .I(N__2003));
    InMux I__211 (
            .O(N__2003),
            .I(N__1999));
    InMux I__210 (
            .O(N__2002),
            .I(N__1996));
    LocalMux I__209 (
            .O(N__1999),
            .I(ctrl_idcodeArea_shifter_3));
    LocalMux I__208 (
            .O(N__1996),
            .I(ctrl_idcodeArea_shifter_3));
    CascadeMux I__207 (
            .O(N__1991),
            .I(N__1987));
    CascadeMux I__206 (
            .O(N__1990),
            .I(N__1984));
    InMux I__205 (
            .O(N__1987),
            .I(N__1979));
    InMux I__204 (
            .O(N__1984),
            .I(N__1979));
    LocalMux I__203 (
            .O(N__1979),
            .I(ctrl_idcodeArea_shifter_2));
    InMux I__202 (
            .O(N__1976),
            .I(N__1970));
    InMux I__201 (
            .O(N__1975),
            .I(N__1970));
    LocalMux I__200 (
            .O(N__1970),
            .I(ctrl_idcodeArea_shifter_7));
    CascadeMux I__199 (
            .O(N__1967),
            .I(N__1963));
    InMux I__198 (
            .O(N__1966),
            .I(N__1958));
    InMux I__197 (
            .O(N__1963),
            .I(N__1958));
    LocalMux I__196 (
            .O(N__1958),
            .I(ctrl_idcodeArea_shifter_10));
    InMux I__195 (
            .O(N__1955),
            .I(N__1949));
    InMux I__194 (
            .O(N__1954),
            .I(N__1949));
    LocalMux I__193 (
            .O(N__1949),
            .I(ctrl_idcodeArea_shifter_9));
    InMux I__192 (
            .O(N__1946),
            .I(N__1940));
    InMux I__191 (
            .O(N__1945),
            .I(N__1940));
    LocalMux I__190 (
            .O(N__1940),
            .I(ctrl_idcodeArea_shifter_8));
    InMux I__189 (
            .O(N__1937),
            .I(N__1931));
    InMux I__188 (
            .O(N__1936),
            .I(N__1931));
    LocalMux I__187 (
            .O(N__1931),
            .I(ctrl_idcodeArea_shifter_4));
    CascadeMux I__186 (
            .O(N__1928),
            .I(N__1925));
    InMux I__185 (
            .O(N__1925),
            .I(N__1919));
    InMux I__184 (
            .O(N__1924),
            .I(N__1919));
    LocalMux I__183 (
            .O(N__1919),
            .I(ctrl_idcodeArea_shifter_6));
    InMux I__182 (
            .O(N__1916),
            .I(N__1910));
    InMux I__181 (
            .O(N__1915),
            .I(N__1910));
    LocalMux I__180 (
            .O(N__1910),
            .I(ctrl_idcodeArea_shifter_5));
    CascadeMux I__179 (
            .O(N__1907),
            .I(N__1903));
    InMux I__178 (
            .O(N__1906),
            .I(N__1900));
    InMux I__177 (
            .O(N__1903),
            .I(N__1897));
    LocalMux I__176 (
            .O(N__1900),
            .I(ctrl_idcodeArea_shifter_11));
    LocalMux I__175 (
            .O(N__1897),
            .I(ctrl_idcodeArea_shifter_11));
    IoInMux I__174 (
            .O(N__1892),
            .I(N__1889));
    LocalMux I__173 (
            .O(N__1889),
            .I(N__1886));
    IoSpan4Mux I__172 (
            .O(N__1886),
            .I(N__1883));
    IoSpan4Mux I__171 (
            .O(N__1883),
            .I(N__1880));
    Span4Mux_s3_h I__170 (
            .O(N__1880),
            .I(N__1876));
    CascadeMux I__169 (
            .O(N__1879),
            .I(N__1873));
    Sp12to4 I__168 (
            .O(N__1876),
            .I(N__1869));
    InMux I__167 (
            .O(N__1873),
            .I(N__1866));
    InMux I__166 (
            .O(N__1872),
            .I(N__1863));
    Odrv12 I__165 (
            .O(N__1869),
            .I(io_leds_c_0));
    LocalMux I__164 (
            .O(N__1866),
            .I(io_leds_c_0));
    LocalMux I__163 (
            .O(N__1863),
            .I(io_leds_c_0));
    IoInMux I__162 (
            .O(N__1856),
            .I(N__1853));
    LocalMux I__161 (
            .O(N__1853),
            .I(N__1850));
    Span4Mux_s3_h I__160 (
            .O(N__1850),
            .I(N__1847));
    Span4Mux_v I__159 (
            .O(N__1847),
            .I(N__1844));
    Sp12to4 I__158 (
            .O(N__1844),
            .I(N__1841));
    Odrv12 I__157 (
            .O(N__1841),
            .I(io_jtag_tck_pad_gb_input));
    defparam IN_MUX_bfv_4_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_7_0_));
    defparam IN_MUX_bfv_4_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_8_0_ (
            .carryinitin(n2066),
            .carryinitout(bfn_4_8_0_));
    defparam IN_MUX_bfv_4_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_9_0_ (
            .carryinitin(n2074),
            .carryinitout(bfn_4_9_0_));
    ICE_GB io_jtag_tck_pad_gb (
            .USERSIGNALTOGLOBALBUFFER(N__1856),
            .GLOBALBUFFEROUTPUT(io_jtag_tck_c));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam ctrl_ledsArea_store_i0_i1_LC_2_5_5.C_ON=1'b0;
    defparam ctrl_ledsArea_store_i0_i1_LC_2_5_5.SEQ_MODE=4'b1000;
    defparam ctrl_ledsArea_store_i0_i1_LC_2_5_5.LUT_INIT=16'b1011101110001000;
    LogicCell40 ctrl_ledsArea_store_i0_i1_LC_2_5_5 (
            .in0(N__1872),
            .in1(N__4415),
            .in2(_gnd_net_),
            .in3(N__2263),
            .lcout(io_leds_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4306),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_ledsArea_shifter_i0_i0_LC_2_6_1.C_ON=1'b0;
    defparam ctrl_ledsArea_shifter_i0_i0_LC_2_6_1.SEQ_MODE=4'b1000;
    defparam ctrl_ledsArea_shifter_i0_i0_LC_2_6_1.LUT_INIT=16'b0011000010101010;
    LogicCell40 ctrl_ledsArea_shifter_i0_i0_LC_2_6_1 (
            .in0(N__4739),
            .in1(N__2093),
            .in2(N__1879),
            .in3(N__4571),
            .lcout(ctrl_ledsArea_shifter_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4305),
            .ce(N__4498),
            .sr(_gnd_net_));
    defparam ctrl_idcodeArea_shifter_i6_LC_4_3_0.C_ON=1'b0;
    defparam ctrl_idcodeArea_shifter_i6_LC_4_3_0.SEQ_MODE=4'b1000;
    defparam ctrl_idcodeArea_shifter_i6_LC_4_3_0.LUT_INIT=16'b1100000010001000;
    LogicCell40 ctrl_idcodeArea_shifter_i6_LC_4_3_0 (
            .in0(N__1975),
            .in1(N__3278),
            .in2(N__1928),
            .in3(N__3423),
            .lcout(ctrl_idcodeArea_shifter_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4316),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_idcodeArea_shifter_i4_LC_4_3_1.C_ON=1'b0;
    defparam ctrl_idcodeArea_shifter_i4_LC_4_3_1.SEQ_MODE=4'b1000;
    defparam ctrl_idcodeArea_shifter_i4_LC_4_3_1.LUT_INIT=16'b1101000010000000;
    LogicCell40 ctrl_idcodeArea_shifter_i4_LC_4_3_1 (
            .in0(N__3421),
            .in1(N__1937),
            .in2(N__3295),
            .in3(N__1915),
            .lcout(ctrl_idcodeArea_shifter_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4316),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_idcodeArea_shifter_i10_LC_4_3_2.C_ON=1'b0;
    defparam ctrl_idcodeArea_shifter_i10_LC_4_3_2.SEQ_MODE=4'b1000;
    defparam ctrl_idcodeArea_shifter_i10_LC_4_3_2.LUT_INIT=16'b1000100011000000;
    LogicCell40 ctrl_idcodeArea_shifter_i10_LC_4_3_2 (
            .in0(N__1966),
            .in1(N__3270),
            .in2(N__1907),
            .in3(N__3419),
            .lcout(ctrl_idcodeArea_shifter_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4316),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_idcodeArea_shifter_i7_LC_4_3_3.C_ON=1'b0;
    defparam ctrl_idcodeArea_shifter_i7_LC_4_3_3.SEQ_MODE=4'b1000;
    defparam ctrl_idcodeArea_shifter_i7_LC_4_3_3.LUT_INIT=16'b1101000010000000;
    LogicCell40 ctrl_idcodeArea_shifter_i7_LC_4_3_3 (
            .in0(N__3424),
            .in1(N__1976),
            .in2(N__3297),
            .in3(N__1945),
            .lcout(ctrl_idcodeArea_shifter_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4316),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_idcodeArea_shifter_i9_LC_4_3_4.C_ON=1'b0;
    defparam ctrl_idcodeArea_shifter_i9_LC_4_3_4.SEQ_MODE=4'b1000;
    defparam ctrl_idcodeArea_shifter_i9_LC_4_3_4.LUT_INIT=16'b1011101111110011;
    LogicCell40 ctrl_idcodeArea_shifter_i9_LC_4_3_4 (
            .in0(N__1955),
            .in1(N__3285),
            .in2(N__1967),
            .in3(N__3426),
            .lcout(ctrl_idcodeArea_shifter_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4316),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_idcodeArea_shifter_i8_LC_4_3_5.C_ON=1'b0;
    defparam ctrl_idcodeArea_shifter_i8_LC_4_3_5.SEQ_MODE=4'b1000;
    defparam ctrl_idcodeArea_shifter_i8_LC_4_3_5.LUT_INIT=16'b1101111110001111;
    LogicCell40 ctrl_idcodeArea_shifter_i8_LC_4_3_5 (
            .in0(N__3425),
            .in1(N__1946),
            .in2(N__3298),
            .in3(N__1954),
            .lcout(ctrl_idcodeArea_shifter_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4316),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_idcodeArea_shifter_i3_LC_4_3_6.C_ON=1'b0;
    defparam ctrl_idcodeArea_shifter_i3_LC_4_3_6.SEQ_MODE=4'b1000;
    defparam ctrl_idcodeArea_shifter_i3_LC_4_3_6.LUT_INIT=16'b1100000010001000;
    LogicCell40 ctrl_idcodeArea_shifter_i3_LC_4_3_6 (
            .in0(N__1936),
            .in1(N__3271),
            .in2(N__2006),
            .in3(N__3420),
            .lcout(ctrl_idcodeArea_shifter_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4316),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_idcodeArea_shifter_i5_LC_4_3_7.C_ON=1'b0;
    defparam ctrl_idcodeArea_shifter_i5_LC_4_3_7.SEQ_MODE=4'b1000;
    defparam ctrl_idcodeArea_shifter_i5_LC_4_3_7.LUT_INIT=16'b1101111110001111;
    LogicCell40 ctrl_idcodeArea_shifter_i5_LC_4_3_7 (
            .in0(N__3422),
            .in1(N__1916),
            .in2(N__3296),
            .in3(N__1924),
            .lcout(ctrl_idcodeArea_shifter_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4316),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_idcodeArea_shifter_i11_LC_4_4_0.C_ON=1'b0;
    defparam ctrl_idcodeArea_shifter_i11_LC_4_4_0.SEQ_MODE=4'b1000;
    defparam ctrl_idcodeArea_shifter_i11_LC_4_4_0.LUT_INIT=16'b1000100011000000;
    LogicCell40 ctrl_idcodeArea_shifter_i11_LC_4_4_0 (
            .in0(N__1906),
            .in1(N__3237),
            .in2(N__2018),
            .in3(N__3401),
            .lcout(ctrl_idcodeArea_shifter_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4312),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_idcodeArea_shifter_i1_LC_4_4_1.C_ON=1'b0;
    defparam ctrl_idcodeArea_shifter_i1_LC_4_4_1.SEQ_MODE=4'b1000;
    defparam ctrl_idcodeArea_shifter_i1_LC_4_4_1.LUT_INIT=16'b1101100000000000;
    LogicCell40 ctrl_idcodeArea_shifter_i1_LC_4_4_1 (
            .in0(N__3407),
            .in1(N__2318),
            .in2(N__1990),
            .in3(N__3243),
            .lcout(ctrl_idcodeArea_shifter_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4312),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_idcodeArea_shifter_i13_LC_4_4_2.C_ON=1'b0;
    defparam ctrl_idcodeArea_shifter_i13_LC_4_4_2.SEQ_MODE=4'b1000;
    defparam ctrl_idcodeArea_shifter_i13_LC_4_4_2.LUT_INIT=16'b1000100011000000;
    LogicCell40 ctrl_idcodeArea_shifter_i13_LC_4_4_2 (
            .in0(N__2029),
            .in1(N__3239),
            .in2(N__2042),
            .in3(N__3403),
            .lcout(ctrl_idcodeArea_shifter_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4312),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_idcodeArea_shifter_i15_LC_4_4_3.C_ON=1'b0;
    defparam ctrl_idcodeArea_shifter_i15_LC_4_4_3.SEQ_MODE=4'b1000;
    defparam ctrl_idcodeArea_shifter_i15_LC_4_4_3.LUT_INIT=16'b1110010000000000;
    LogicCell40 ctrl_idcodeArea_shifter_i15_LC_4_4_3 (
            .in0(N__3405),
            .in1(N__2065),
            .in2(N__2057),
            .in3(N__3242),
            .lcout(ctrl_idcodeArea_shifter_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4312),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_idcodeArea_shifter_i16_LC_4_4_4.C_ON=1'b0;
    defparam ctrl_idcodeArea_shifter_i16_LC_4_4_4.SEQ_MODE=4'b1000;
    defparam ctrl_idcodeArea_shifter_i16_LC_4_4_4.LUT_INIT=16'b1011101111110011;
    LogicCell40 ctrl_idcodeArea_shifter_i16_LC_4_4_4 (
            .in0(N__2066),
            .in1(N__3240),
            .in2(N__2336),
            .in3(N__3406),
            .lcout(ctrl_idcodeArea_shifter_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4312),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_idcodeArea_shifter_i14_LC_4_4_5.C_ON=1'b0;
    defparam ctrl_idcodeArea_shifter_i14_LC_4_4_5.SEQ_MODE=4'b1000;
    defparam ctrl_idcodeArea_shifter_i14_LC_4_4_5.LUT_INIT=16'b1101100011111111;
    LogicCell40 ctrl_idcodeArea_shifter_i14_LC_4_4_5 (
            .in0(N__3404),
            .in1(N__2041),
            .in2(N__2056),
            .in3(N__3241),
            .lcout(ctrl_idcodeArea_shifter_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4312),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_idcodeArea_shifter_i12_LC_4_4_6.C_ON=1'b0;
    defparam ctrl_idcodeArea_shifter_i12_LC_4_4_6.SEQ_MODE=4'b1000;
    defparam ctrl_idcodeArea_shifter_i12_LC_4_4_6.LUT_INIT=16'b1000100011000000;
    LogicCell40 ctrl_idcodeArea_shifter_i12_LC_4_4_6 (
            .in0(N__2017),
            .in1(N__3238),
            .in2(N__2030),
            .in3(N__3402),
            .lcout(ctrl_idcodeArea_shifter_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4312),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_idcodeArea_shifter_i2_LC_4_4_7.C_ON=1'b0;
    defparam ctrl_idcodeArea_shifter_i2_LC_4_4_7.SEQ_MODE=4'b1000;
    defparam ctrl_idcodeArea_shifter_i2_LC_4_4_7.LUT_INIT=16'b1110010000000000;
    LogicCell40 ctrl_idcodeArea_shifter_i2_LC_4_4_7 (
            .in0(N__3408),
            .in1(N__2002),
            .in2(N__1991),
            .in3(N__3244),
            .lcout(ctrl_idcodeArea_shifter_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4312),
            .ce(),
            .sr(_gnd_net_));
    defparam i1546_2_lut_3_lut_LC_4_5_0.C_ON=1'b0;
    defparam i1546_2_lut_3_lut_LC_4_5_0.SEQ_MODE=4'b0000;
    defparam i1546_2_lut_3_lut_LC_4_5_0.LUT_INIT=16'b1100110011101110;
    LogicCell40 i1546_2_lut_3_lut_LC_4_5_0 (
            .in0(N__3819),
            .in1(N__3912),
            .in2(_gnd_net_),
            .in3(N__3721),
            .lcout(n2248),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1457_2_lut_LC_4_5_1.C_ON=1'b0;
    defparam i1457_2_lut_LC_4_5_1.SEQ_MODE=4'b0000;
    defparam i1457_2_lut_LC_4_5_1.LUT_INIT=16'b1100110000000000;
    LogicCell40 i1457_2_lut_LC_4_5_1 (
            .in0(_gnd_net_),
            .in1(N__3703),
            .in2(_gnd_net_),
            .in3(N__3818),
            .lcout(n2206),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1555_2_lut_LC_4_5_2.C_ON=1'b0;
    defparam i1555_2_lut_LC_4_5_2.SEQ_MODE=4'b0000;
    defparam i1555_2_lut_LC_4_5_2.LUT_INIT=16'b1111111100110011;
    LogicCell40 i1555_2_lut_LC_4_5_2 (
            .in0(_gnd_net_),
            .in1(N__4199),
            .in2(_gnd_net_),
            .in3(N__3722),
            .lcout(n2306),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_tap_instructionShift_i0_i0_LC_4_5_3.C_ON=1'b0;
    defparam ctrl_tap_instructionShift_i0_i0_LC_4_5_3.SEQ_MODE=4'b1000;
    defparam ctrl_tap_instructionShift_i0_i0_LC_4_5_3.LUT_INIT=16'b1100110010101010;
    LogicCell40 ctrl_tap_instructionShift_i0_i0_LC_4_5_3 (
            .in0(N__2389),
            .in1(N__2521),
            .in2(_gnd_net_),
            .in3(N__3704),
            .lcout(ctrl_tap_instructionShift_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4309),
            .ce(N__2566),
            .sr(_gnd_net_));
    defparam ctrl_tap_instructionShift_i0_i1_LC_4_5_4.C_ON=1'b0;
    defparam ctrl_tap_instructionShift_i0_i1_LC_4_5_4.SEQ_MODE=4'b1000;
    defparam ctrl_tap_instructionShift_i0_i1_LC_4_5_4.LUT_INIT=16'b1100110010101010;
    LogicCell40 ctrl_tap_instructionShift_i0_i1_LC_4_5_4 (
            .in0(N__2443),
            .in1(N__2377),
            .in2(_gnd_net_),
            .in3(N__3723),
            .lcout(ctrl_tap_instructionShift_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4309),
            .ce(N__2566),
            .sr(_gnd_net_));
    defparam ctrl_tap_instructionShift_i0_i2_LC_4_5_5.C_ON=1'b0;
    defparam ctrl_tap_instructionShift_i0_i2_LC_4_5_5.SEQ_MODE=4'b1000;
    defparam ctrl_tap_instructionShift_i0_i2_LC_4_5_5.LUT_INIT=16'b1100110010101010;
    LogicCell40 ctrl_tap_instructionShift_i0_i2_LC_4_5_5 (
            .in0(N__2491),
            .in1(N__2431),
            .in2(_gnd_net_),
            .in3(N__3705),
            .lcout(ctrl_tap_instructionShift_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4309),
            .ce(N__2566),
            .sr(_gnd_net_));
    defparam ctrl_tap_instructionShift_i0_i3_LC_4_5_6.C_ON=1'b0;
    defparam ctrl_tap_instructionShift_i0_i3_LC_4_5_6.SEQ_MODE=4'b1000;
    defparam ctrl_tap_instructionShift_i0_i3_LC_4_5_6.LUT_INIT=16'b1100110010101010;
    LogicCell40 ctrl_tap_instructionShift_i0_i3_LC_4_5_6 (
            .in0(N__3522),
            .in1(N__2480),
            .in2(_gnd_net_),
            .in3(N__3724),
            .lcout(ctrl_tap_instructionShift_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4309),
            .ce(N__2566),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_4_lut_adj_2_LC_4_6_2.C_ON=1'b0;
    defparam i1_2_lut_3_lut_4_lut_adj_2_LC_4_6_2.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_4_lut_adj_2_LC_4_6_2.LUT_INIT=16'b1110111111111111;
    LogicCell40 i1_2_lut_3_lut_4_lut_adj_2_LC_4_6_2 (
            .in0(N__3715),
            .in1(N__4034),
            .in2(N__4160),
            .in3(N__3837),
            .lcout(n7),
            .ltout(n7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_ledsArea_shifter_i0_i7_LC_4_6_3.C_ON=1'b0;
    defparam ctrl_ledsArea_shifter_i0_i7_LC_4_6_3.SEQ_MODE=4'b1000;
    defparam ctrl_ledsArea_shifter_i0_i7_LC_4_6_3.LUT_INIT=16'b0000110010101010;
    LogicCell40 ctrl_ledsArea_shifter_i0_i7_LC_4_6_3 (
            .in0(N__3524),
            .in1(N__2796),
            .in2(N__2084),
            .in3(N__4570),
            .lcout(ctrl_ledsArea_shifter_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4307),
            .ce(N__4497),
            .sr(_gnd_net_));
    defparam i1_2_lut_4_lut_LC_4_6_5.C_ON=1'b0;
    defparam i1_2_lut_4_lut_LC_4_6_5.SEQ_MODE=4'b0000;
    defparam i1_2_lut_4_lut_LC_4_6_5.LUT_INIT=16'b0000000000001000;
    LogicCell40 i1_2_lut_4_lut_LC_4_6_5 (
            .in0(N__3836),
            .in1(N__4156),
            .in2(N__2285),
            .in3(N__4035),
            .lcout(n1275),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_4_lut_LC_4_6_6.C_ON=1'b0;
    defparam i1_2_lut_3_lut_4_lut_LC_4_6_6.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_4_lut_LC_4_6_6.LUT_INIT=16'b1101111111111111;
    LogicCell40 i1_2_lut_3_lut_4_lut_LC_4_6_6 (
            .in0(N__2520),
            .in1(N__2474),
            .in2(N__2378),
            .in3(N__2430),
            .lcout(n7_adj_1),
            .ltout(n7_adj_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i4_4_lut_LC_4_6_7.C_ON=1'b0;
    defparam i4_4_lut_LC_4_6_7.SEQ_MODE=4'b0000;
    defparam i4_4_lut_LC_4_6_7.LUT_INIT=16'b1111011111111111;
    LogicCell40 i4_4_lut_LC_4_6_7 (
            .in0(N__4033),
            .in1(N__2081),
            .in2(N__2075),
            .in3(N__4155),
            .lcout(n2110),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam myClockArea_timeout_counter_value_317__i0_LC_4_7_0.C_ON=1'b1;
    defparam myClockArea_timeout_counter_value_317__i0_LC_4_7_0.SEQ_MODE=4'b1010;
    defparam myClockArea_timeout_counter_value_317__i0_LC_4_7_0.LUT_INIT=16'b1000001000101000;
    LogicCell40 myClockArea_timeout_counter_value_317__i0_LC_4_7_0 (
            .in0(N__3108),
            .in1(N__2738),
            .in2(_gnd_net_),
            .in3(N__2072),
            .lcout(myClockArea_timeout_counter_value_0),
            .ltout(),
            .carryin(bfn_4_7_0_),
            .carryout(n2059),
            .clk(N__2846),
            .ce(),
            .sr(N__2227));
    defparam myClockArea_timeout_counter_value_317__i1_LC_4_7_1.C_ON=1'b1;
    defparam myClockArea_timeout_counter_value_317__i1_LC_4_7_1.SEQ_MODE=4'b1010;
    defparam myClockArea_timeout_counter_value_317__i1_LC_4_7_1.LUT_INIT=16'b1000001000101000;
    LogicCell40 myClockArea_timeout_counter_value_317__i1_LC_4_7_1 (
            .in0(N__3095),
            .in1(N__2765),
            .in2(_gnd_net_),
            .in3(N__2069),
            .lcout(myClockArea_timeout_counter_value_1),
            .ltout(),
            .carryin(n2059),
            .carryout(n2060),
            .clk(N__2846),
            .ce(),
            .sr(N__2227));
    defparam myClockArea_timeout_counter_value_317__i2_LC_4_7_2.C_ON=1'b1;
    defparam myClockArea_timeout_counter_value_317__i2_LC_4_7_2.SEQ_MODE=4'b1010;
    defparam myClockArea_timeout_counter_value_317__i2_LC_4_7_2.LUT_INIT=16'b1000001000101000;
    LogicCell40 myClockArea_timeout_counter_value_317__i2_LC_4_7_2 (
            .in0(N__3109),
            .in1(N__2630),
            .in2(_gnd_net_),
            .in3(N__2120),
            .lcout(myClockArea_timeout_counter_value_2),
            .ltout(),
            .carryin(n2060),
            .carryout(n2061),
            .clk(N__2846),
            .ce(),
            .sr(N__2227));
    defparam myClockArea_timeout_counter_value_317__i3_LC_4_7_3.C_ON=1'b1;
    defparam myClockArea_timeout_counter_value_317__i3_LC_4_7_3.SEQ_MODE=4'b1010;
    defparam myClockArea_timeout_counter_value_317__i3_LC_4_7_3.LUT_INIT=16'b1000001000101000;
    LogicCell40 myClockArea_timeout_counter_value_317__i3_LC_4_7_3 (
            .in0(N__3096),
            .in1(N__2777),
            .in2(_gnd_net_),
            .in3(N__2117),
            .lcout(myClockArea_timeout_counter_value_3),
            .ltout(),
            .carryin(n2061),
            .carryout(n2062),
            .clk(N__2846),
            .ce(),
            .sr(N__2227));
    defparam myClockArea_timeout_counter_value_317__i4_LC_4_7_4.C_ON=1'b1;
    defparam myClockArea_timeout_counter_value_317__i4_LC_4_7_4.SEQ_MODE=4'b1010;
    defparam myClockArea_timeout_counter_value_317__i4_LC_4_7_4.LUT_INIT=16'b1000001000101000;
    LogicCell40 myClockArea_timeout_counter_value_317__i4_LC_4_7_4 (
            .in0(N__3110),
            .in1(N__2720),
            .in2(_gnd_net_),
            .in3(N__2114),
            .lcout(myClockArea_timeout_counter_value_4),
            .ltout(),
            .carryin(n2062),
            .carryout(n2063),
            .clk(N__2846),
            .ce(),
            .sr(N__2227));
    defparam myClockArea_timeout_counter_value_317__i5_LC_4_7_5.C_ON=1'b1;
    defparam myClockArea_timeout_counter_value_317__i5_LC_4_7_5.SEQ_MODE=4'b1010;
    defparam myClockArea_timeout_counter_value_317__i5_LC_4_7_5.LUT_INIT=16'b1000001000101000;
    LogicCell40 myClockArea_timeout_counter_value_317__i5_LC_4_7_5 (
            .in0(N__3097),
            .in1(N__2752),
            .in2(_gnd_net_),
            .in3(N__2111),
            .lcout(myClockArea_timeout_counter_value_5),
            .ltout(),
            .carryin(n2063),
            .carryout(n2064),
            .clk(N__2846),
            .ce(),
            .sr(N__2227));
    defparam myClockArea_timeout_counter_value_317__i6_LC_4_7_6.C_ON=1'b1;
    defparam myClockArea_timeout_counter_value_317__i6_LC_4_7_6.SEQ_MODE=4'b1010;
    defparam myClockArea_timeout_counter_value_317__i6_LC_4_7_6.LUT_INIT=16'b1000001000101000;
    LogicCell40 myClockArea_timeout_counter_value_317__i6_LC_4_7_6 (
            .in0(N__3111),
            .in1(N__2708),
            .in2(_gnd_net_),
            .in3(N__2108),
            .lcout(myClockArea_timeout_counter_value_6),
            .ltout(),
            .carryin(n2064),
            .carryout(n2065),
            .clk(N__2846),
            .ce(),
            .sr(N__2227));
    defparam myClockArea_timeout_counter_value_317__i7_LC_4_7_7.C_ON=1'b1;
    defparam myClockArea_timeout_counter_value_317__i7_LC_4_7_7.SEQ_MODE=4'b1010;
    defparam myClockArea_timeout_counter_value_317__i7_LC_4_7_7.LUT_INIT=16'b1000001000101000;
    LogicCell40 myClockArea_timeout_counter_value_317__i7_LC_4_7_7 (
            .in0(N__3098),
            .in1(N__3029),
            .in2(_gnd_net_),
            .in3(N__2105),
            .lcout(myClockArea_timeout_counter_value_7),
            .ltout(),
            .carryin(n2065),
            .carryout(n2066),
            .clk(N__2846),
            .ce(),
            .sr(N__2227));
    defparam myClockArea_timeout_counter_value_317__i8_LC_4_8_0.C_ON=1'b1;
    defparam myClockArea_timeout_counter_value_317__i8_LC_4_8_0.SEQ_MODE=4'b1010;
    defparam myClockArea_timeout_counter_value_317__i8_LC_4_8_0.LUT_INIT=16'b1000001000101000;
    LogicCell40 myClockArea_timeout_counter_value_317__i8_LC_4_8_0 (
            .in0(N__3119),
            .in1(N__2657),
            .in2(_gnd_net_),
            .in3(N__2102),
            .lcout(myClockArea_timeout_counter_value_8),
            .ltout(),
            .carryin(bfn_4_8_0_),
            .carryout(n2067),
            .clk(N__2845),
            .ce(),
            .sr(N__2228));
    defparam myClockArea_timeout_counter_value_317__i9_LC_4_8_1.C_ON=1'b1;
    defparam myClockArea_timeout_counter_value_317__i9_LC_4_8_1.SEQ_MODE=4'b1010;
    defparam myClockArea_timeout_counter_value_317__i9_LC_4_8_1.LUT_INIT=16'b1000001000101000;
    LogicCell40 myClockArea_timeout_counter_value_317__i9_LC_4_8_1 (
            .in0(N__3091),
            .in1(N__2942),
            .in2(_gnd_net_),
            .in3(N__2099),
            .lcout(myClockArea_timeout_counter_value_9),
            .ltout(),
            .carryin(n2067),
            .carryout(n2068),
            .clk(N__2845),
            .ce(),
            .sr(N__2228));
    defparam myClockArea_timeout_counter_value_317__i10_LC_4_8_2.C_ON=1'b1;
    defparam myClockArea_timeout_counter_value_317__i10_LC_4_8_2.SEQ_MODE=4'b1010;
    defparam myClockArea_timeout_counter_value_317__i10_LC_4_8_2.LUT_INIT=16'b1000001000101000;
    LogicCell40 myClockArea_timeout_counter_value_317__i10_LC_4_8_2 (
            .in0(N__3116),
            .in1(N__2644),
            .in2(_gnd_net_),
            .in3(N__2096),
            .lcout(myClockArea_timeout_counter_value_10),
            .ltout(),
            .carryin(n2068),
            .carryout(n2069),
            .clk(N__2845),
            .ce(),
            .sr(N__2228));
    defparam myClockArea_timeout_counter_value_317__i11_LC_4_8_3.C_ON=1'b1;
    defparam myClockArea_timeout_counter_value_317__i11_LC_4_8_3.SEQ_MODE=4'b1010;
    defparam myClockArea_timeout_counter_value_317__i11_LC_4_8_3.LUT_INIT=16'b1000001000101000;
    LogicCell40 myClockArea_timeout_counter_value_317__i11_LC_4_8_3 (
            .in0(N__3088),
            .in1(N__2960),
            .in2(_gnd_net_),
            .in3(N__2147),
            .lcout(myClockArea_timeout_counter_value_11),
            .ltout(),
            .carryin(n2069),
            .carryout(n2070),
            .clk(N__2845),
            .ce(),
            .sr(N__2228));
    defparam myClockArea_timeout_counter_value_317__i12_LC_4_8_4.C_ON=1'b1;
    defparam myClockArea_timeout_counter_value_317__i12_LC_4_8_4.SEQ_MODE=4'b1010;
    defparam myClockArea_timeout_counter_value_317__i12_LC_4_8_4.LUT_INIT=16'b1000001000101000;
    LogicCell40 myClockArea_timeout_counter_value_317__i12_LC_4_8_4 (
            .in0(N__3117),
            .in1(N__2917),
            .in2(_gnd_net_),
            .in3(N__2144),
            .lcout(myClockArea_timeout_counter_value_12),
            .ltout(),
            .carryin(n2070),
            .carryout(n2071),
            .clk(N__2845),
            .ce(),
            .sr(N__2228));
    defparam myClockArea_timeout_counter_value_317__i13_LC_4_8_5.C_ON=1'b1;
    defparam myClockArea_timeout_counter_value_317__i13_LC_4_8_5.SEQ_MODE=4'b1010;
    defparam myClockArea_timeout_counter_value_317__i13_LC_4_8_5.LUT_INIT=16'b1000001000101000;
    LogicCell40 myClockArea_timeout_counter_value_317__i13_LC_4_8_5 (
            .in0(N__3089),
            .in1(N__2603),
            .in2(_gnd_net_),
            .in3(N__2141),
            .lcout(myClockArea_timeout_counter_value_13),
            .ltout(),
            .carryin(n2071),
            .carryout(n2072),
            .clk(N__2845),
            .ce(),
            .sr(N__2228));
    defparam myClockArea_timeout_counter_value_317__i14_LC_4_8_6.C_ON=1'b1;
    defparam myClockArea_timeout_counter_value_317__i14_LC_4_8_6.SEQ_MODE=4'b1010;
    defparam myClockArea_timeout_counter_value_317__i14_LC_4_8_6.LUT_INIT=16'b1000001000101000;
    LogicCell40 myClockArea_timeout_counter_value_317__i14_LC_4_8_6 (
            .in0(N__3118),
            .in1(N__2903),
            .in2(_gnd_net_),
            .in3(N__2138),
            .lcout(myClockArea_timeout_counter_value_14),
            .ltout(),
            .carryin(n2072),
            .carryout(n2073),
            .clk(N__2845),
            .ce(),
            .sr(N__2228));
    defparam myClockArea_timeout_counter_value_317__i15_LC_4_8_7.C_ON=1'b1;
    defparam myClockArea_timeout_counter_value_317__i15_LC_4_8_7.SEQ_MODE=4'b1010;
    defparam myClockArea_timeout_counter_value_317__i15_LC_4_8_7.LUT_INIT=16'b1000001000101000;
    LogicCell40 myClockArea_timeout_counter_value_317__i15_LC_4_8_7 (
            .in0(N__3090),
            .in1(N__2987),
            .in2(_gnd_net_),
            .in3(N__2135),
            .lcout(myClockArea_timeout_counter_value_15),
            .ltout(),
            .carryin(n2073),
            .carryout(n2074),
            .clk(N__2845),
            .ce(),
            .sr(N__2228));
    defparam myClockArea_timeout_counter_value_317__i16_LC_4_9_0.C_ON=1'b1;
    defparam myClockArea_timeout_counter_value_317__i16_LC_4_9_0.SEQ_MODE=4'b1010;
    defparam myClockArea_timeout_counter_value_317__i16_LC_4_9_0.LUT_INIT=16'b1000001000101000;
    LogicCell40 myClockArea_timeout_counter_value_317__i16_LC_4_9_0 (
            .in0(N__3112),
            .in1(N__2681),
            .in2(_gnd_net_),
            .in3(N__2132),
            .lcout(myClockArea_timeout_counter_value_16),
            .ltout(),
            .carryin(bfn_4_9_0_),
            .carryout(n2075),
            .clk(N__2847),
            .ce(),
            .sr(N__2223));
    defparam myClockArea_timeout_counter_value_317__i17_LC_4_9_1.C_ON=1'b1;
    defparam myClockArea_timeout_counter_value_317__i17_LC_4_9_1.SEQ_MODE=4'b1010;
    defparam myClockArea_timeout_counter_value_317__i17_LC_4_9_1.LUT_INIT=16'b1000001000101000;
    LogicCell40 myClockArea_timeout_counter_value_317__i17_LC_4_9_1 (
            .in0(N__3092),
            .in1(N__2669),
            .in2(_gnd_net_),
            .in3(N__2129),
            .lcout(myClockArea_timeout_counter_value_17),
            .ltout(),
            .carryin(n2075),
            .carryout(n2076),
            .clk(N__2847),
            .ce(),
            .sr(N__2223));
    defparam myClockArea_timeout_counter_value_317__i18_LC_4_9_2.C_ON=1'b1;
    defparam myClockArea_timeout_counter_value_317__i18_LC_4_9_2.SEQ_MODE=4'b1010;
    defparam myClockArea_timeout_counter_value_317__i18_LC_4_9_2.LUT_INIT=16'b1000001000101000;
    LogicCell40 myClockArea_timeout_counter_value_317__i18_LC_4_9_2 (
            .in0(N__3113),
            .in1(N__2930),
            .in2(_gnd_net_),
            .in3(N__2126),
            .lcout(myClockArea_timeout_counter_value_18),
            .ltout(),
            .carryin(n2076),
            .carryout(n2077),
            .clk(N__2847),
            .ce(),
            .sr(N__2223));
    defparam myClockArea_timeout_counter_value_317__i19_LC_4_9_3.C_ON=1'b1;
    defparam myClockArea_timeout_counter_value_317__i19_LC_4_9_3.SEQ_MODE=4'b1010;
    defparam myClockArea_timeout_counter_value_317__i19_LC_4_9_3.LUT_INIT=16'b1000001000101000;
    LogicCell40 myClockArea_timeout_counter_value_317__i19_LC_4_9_3 (
            .in0(N__3093),
            .in1(N__2999),
            .in2(_gnd_net_),
            .in3(N__2123),
            .lcout(myClockArea_timeout_counter_value_19),
            .ltout(),
            .carryin(n2077),
            .carryout(n2078),
            .clk(N__2847),
            .ce(),
            .sr(N__2223));
    defparam myClockArea_timeout_counter_value_317__i20_LC_4_9_4.C_ON=1'b1;
    defparam myClockArea_timeout_counter_value_317__i20_LC_4_9_4.SEQ_MODE=4'b1010;
    defparam myClockArea_timeout_counter_value_317__i20_LC_4_9_4.LUT_INIT=16'b1000001000101000;
    LogicCell40 myClockArea_timeout_counter_value_317__i20_LC_4_9_4 (
            .in0(N__3114),
            .in1(N__2974),
            .in2(_gnd_net_),
            .in3(N__2237),
            .lcout(myClockArea_timeout_counter_value_20),
            .ltout(),
            .carryin(n2078),
            .carryout(n2079),
            .clk(N__2847),
            .ce(),
            .sr(N__2223));
    defparam myClockArea_timeout_counter_value_317__i21_LC_4_9_5.C_ON=1'b1;
    defparam myClockArea_timeout_counter_value_317__i21_LC_4_9_5.SEQ_MODE=4'b1010;
    defparam myClockArea_timeout_counter_value_317__i21_LC_4_9_5.LUT_INIT=16'b1000001000101000;
    LogicCell40 myClockArea_timeout_counter_value_317__i21_LC_4_9_5 (
            .in0(N__3094),
            .in1(N__3017),
            .in2(_gnd_net_),
            .in3(N__2234),
            .lcout(myClockArea_timeout_counter_value_21),
            .ltout(),
            .carryin(n2079),
            .carryout(n2080),
            .clk(N__2847),
            .ce(),
            .sr(N__2223));
    defparam myClockArea_timeout_counter_value_317__i22_LC_4_9_6.C_ON=1'b0;
    defparam myClockArea_timeout_counter_value_317__i22_LC_4_9_6.SEQ_MODE=4'b1010;
    defparam myClockArea_timeout_counter_value_317__i22_LC_4_9_6.LUT_INIT=16'b1000001000101000;
    LogicCell40 myClockArea_timeout_counter_value_317__i22_LC_4_9_6 (
            .in0(N__3115),
            .in1(N__2695),
            .in2(_gnd_net_),
            .in3(N__2231),
            .lcout(myClockArea_timeout_counter_value_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2847),
            .ce(),
            .sr(N__2223));
    defparam myClockArea_timeout_state_90_LC_4_10_0.C_ON=1'b0;
    defparam myClockArea_timeout_state_90_LC_4_10_0.SEQ_MODE=4'b1010;
    defparam myClockArea_timeout_state_90_LC_4_10_0.LUT_INIT=16'b0000000001010101;
    LogicCell40 myClockArea_timeout_state_90_LC_4_10_0 (
            .in0(N__2588),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2883),
            .lcout(myClockArea_timeout_state),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2848),
            .ce(),
            .sr(N__2213));
    defparam ctrl_idcodeArea_shifter_i28_LC_5_3_2.C_ON=1'b0;
    defparam ctrl_idcodeArea_shifter_i28_LC_5_3_2.SEQ_MODE=4'b1000;
    defparam ctrl_idcodeArea_shifter_i28_LC_5_3_2.LUT_INIT=16'b1101000010000000;
    LogicCell40 ctrl_idcodeArea_shifter_i28_LC_5_3_2 (
            .in0(N__3415),
            .in1(N__2177),
            .in2(N__3292),
            .in3(N__2155),
            .lcout(ctrl_idcodeArea_shifter_28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4319),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_idcodeArea_shifter_i30_LC_5_3_3.C_ON=1'b0;
    defparam ctrl_idcodeArea_shifter_i30_LC_5_3_3.SEQ_MODE=4'b1000;
    defparam ctrl_idcodeArea_shifter_i30_LC_5_3_3.LUT_INIT=16'b1100000010001000;
    LogicCell40 ctrl_idcodeArea_shifter_i30_LC_5_3_3 (
            .in0(N__2185),
            .in1(N__3266),
            .in2(N__2168),
            .in3(N__3417),
            .lcout(ctrl_idcodeArea_shifter_30),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4319),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_idcodeArea_shifter_i31_LC_5_3_4.C_ON=1'b0;
    defparam ctrl_idcodeArea_shifter_i31_LC_5_3_4.SEQ_MODE=4'b1000;
    defparam ctrl_idcodeArea_shifter_i31_LC_5_3_4.LUT_INIT=16'b1110111101001111;
    LogicCell40 ctrl_idcodeArea_shifter_i31_LC_5_3_4 (
            .in0(N__3418),
            .in1(N__3512),
            .in2(N__3294),
            .in3(N__2186),
            .lcout(ctrl_idcodeArea_shifter_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4319),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_idcodeArea_shifter_i27_LC_5_3_5.C_ON=1'b0;
    defparam ctrl_idcodeArea_shifter_i27_LC_5_3_5.SEQ_MODE=4'b1000;
    defparam ctrl_idcodeArea_shifter_i27_LC_5_3_5.LUT_INIT=16'b1100000010001000;
    LogicCell40 ctrl_idcodeArea_shifter_i27_LC_5_3_5 (
            .in0(N__2176),
            .in1(N__3259),
            .in2(N__3554),
            .in3(N__3414),
            .lcout(ctrl_idcodeArea_shifter_27),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4319),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_idcodeArea_shifter_i29_LC_5_3_6.C_ON=1'b0;
    defparam ctrl_idcodeArea_shifter_i29_LC_5_3_6.SEQ_MODE=4'b1000;
    defparam ctrl_idcodeArea_shifter_i29_LC_5_3_6.LUT_INIT=16'b1101000010000000;
    LogicCell40 ctrl_idcodeArea_shifter_i29_LC_5_3_6 (
            .in0(N__3416),
            .in1(N__2156),
            .in2(N__3293),
            .in3(N__2164),
            .lcout(ctrl_idcodeArea_shifter_29),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4319),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_idcodeArea_shifter_i17_LC_5_4_0.C_ON=1'b0;
    defparam ctrl_idcodeArea_shifter_i17_LC_5_4_0.SEQ_MODE=4'b1000;
    defparam ctrl_idcodeArea_shifter_i17_LC_5_4_0.LUT_INIT=16'b1101100000000000;
    LogicCell40 ctrl_idcodeArea_shifter_i17_LC_5_4_0 (
            .in0(N__3400),
            .in1(N__2332),
            .in2(N__3446),
            .in3(N__3208),
            .lcout(ctrl_idcodeArea_shifter_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4317),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_3_lut_4_lut_adj_5_LC_5_4_1.C_ON=1'b0;
    defparam i2_3_lut_4_lut_adj_5_LC_5_4_1.SEQ_MODE=4'b0000;
    defparam i2_3_lut_4_lut_adj_5_LC_5_4_1.LUT_INIT=16'b1111101111111111;
    LogicCell40 i2_3_lut_4_lut_adj_5_LC_5_4_1 (
            .in0(N__2428),
            .in1(N__2372),
            .in2(N__2479),
            .in3(N__2518),
            .lcout(n2085),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_idcodeArea_shifter_i0_LC_5_4_2.C_ON=1'b0;
    defparam ctrl_idcodeArea_shifter_i0_LC_5_4_2.SEQ_MODE=4'b1000;
    defparam ctrl_idcodeArea_shifter_i0_LC_5_4_2.LUT_INIT=16'b1010110011111111;
    LogicCell40 ctrl_idcodeArea_shifter_i0_LC_5_4_2 (
            .in0(N__2303),
            .in1(N__2317),
            .in2(N__3431),
            .in3(N__3207),
            .lcout(ctrl_idcodeArea_shifter_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4317),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_ledsArea_store_i0_i6_LC_5_4_3.C_ON=1'b0;
    defparam ctrl_ledsArea_store_i0_i6_LC_5_4_3.SEQ_MODE=4'b1000;
    defparam ctrl_ledsArea_store_i0_i6_LC_5_4_3.LUT_INIT=16'b1100110010101010;
    LogicCell40 ctrl_ledsArea_store_i0_i6_LC_5_4_3 (
            .in0(N__4664),
            .in1(N__4677),
            .in2(_gnd_net_),
            .in3(N__4418),
            .lcout(io_leds_c_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4317),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_tap_instruction_3__I_0_i6_2_lut_LC_5_4_4.C_ON=1'b0;
    defparam ctrl_tap_instruction_3__I_0_i6_2_lut_LC_5_4_4.SEQ_MODE=4'b0000;
    defparam ctrl_tap_instruction_3__I_0_i6_2_lut_LC_5_4_4.LUT_INIT=16'b1111111100110011;
    LogicCell40 ctrl_tap_instruction_3__I_0_i6_2_lut_LC_5_4_4 (
            .in0(_gnd_net_),
            .in1(N__2429),
            .in2(_gnd_net_),
            .in3(N__2470),
            .lcout(),
            .ltout(n6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam equal_316_i15_4_lut_LC_5_4_5.C_ON=1'b0;
    defparam equal_316_i15_4_lut_LC_5_4_5.SEQ_MODE=4'b0000;
    defparam equal_316_i15_4_lut_LC_5_4_5.LUT_INIT=16'b1111111111111110;
    LogicCell40 equal_316_i15_4_lut_LC_5_4_5 (
            .in0(N__2371),
            .in1(N__2519),
            .in2(N__2306),
            .in3(N__4551),
            .lcout(n15),
            .ltout(n15_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i397_4_lut_LC_5_4_6.C_ON=1'b0;
    defparam i397_4_lut_LC_5_4_6.SEQ_MODE=4'b0000;
    defparam i397_4_lut_LC_5_4_6.LUT_INIT=16'b1100101000001010;
    LogicCell40 i397_4_lut_LC_5_4_6 (
            .in0(N__2302),
            .in1(N__2294),
            .in2(N__2288),
            .in3(N__3560),
            .lcout(),
            .ltout(ctrl_tap_tdoUnbufferd_N_211_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i400_4_lut_LC_5_4_7.C_ON=1'b0;
    defparam i400_4_lut_LC_5_4_7.SEQ_MODE=4'b0000;
    defparam i400_4_lut_LC_5_4_7.LUT_INIT=16'b1111000011100100;
    LogicCell40 i400_4_lut_LC_5_4_7 (
            .in0(N__2284),
            .in1(N__2267),
            .in2(N__2249),
            .in3(N__4552),
            .lcout(ctrl_tap_tdoUnbufferd),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_3_lut_4_lut_adj_3_LC_5_5_0.C_ON=1'b0;
    defparam i2_3_lut_4_lut_adj_3_LC_5_5_0.SEQ_MODE=4'b0000;
    defparam i2_3_lut_4_lut_adj_3_LC_5_5_0.LUT_INIT=16'b1111111111111110;
    LogicCell40 i2_3_lut_4_lut_adj_3_LC_5_5_0 (
            .in0(N__3838),
            .in1(N__3711),
            .in2(N__4154),
            .in3(N__4039),
            .lcout(n1489),
            .ltout(n1489_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_4_lut_LC_5_5_1.C_ON=1'b0;
    defparam i1_3_lut_4_lut_LC_5_5_1.SEQ_MODE=4'b0000;
    defparam i1_3_lut_4_lut_LC_5_5_1.LUT_INIT=16'b0001111100001111;
    LogicCell40 i1_3_lut_4_lut_LC_5_5_1 (
            .in0(N__4040),
            .in1(N__3596),
            .in2(N__2528),
            .in3(N__4141),
            .lcout(n1269),
            .ltout(n1269_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_tap_instruction_i0_LC_5_5_2.C_ON=1'b0;
    defparam ctrl_tap_instruction_i0_LC_5_5_2.SEQ_MODE=4'b1000;
    defparam ctrl_tap_instruction_i0_LC_5_5_2.LUT_INIT=16'b1010110000001100;
    LogicCell40 ctrl_tap_instruction_i0_LC_5_5_2 (
            .in0(N__3206),
            .in1(N__2522),
            .in2(N__2525),
            .in3(N__3589),
            .lcout(ctrl_tap_instruction_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4313),
            .ce(),
            .sr(_gnd_net_));
    defparam i917_4_lut_4_lut_LC_5_5_3.C_ON=1'b0;
    defparam i917_4_lut_4_lut_LC_5_5_3.SEQ_MODE=4'b0000;
    defparam i917_4_lut_4_lut_LC_5_5_3.LUT_INIT=16'b0001000000000010;
    LogicCell40 i917_4_lut_4_lut_LC_5_5_3 (
            .in0(N__4038),
            .in1(N__4140),
            .in2(N__3732),
            .in3(N__3839),
            .lcout(n1022),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_tap_instruction_i3_LC_5_5_4.C_ON=1'b0;
    defparam ctrl_tap_instruction_i3_LC_5_5_4.SEQ_MODE=4'b1000;
    defparam ctrl_tap_instruction_i3_LC_5_5_4.LUT_INIT=16'b1010001010000000;
    LogicCell40 ctrl_tap_instruction_i3_LC_5_5_4 (
            .in0(N__3205),
            .in1(N__2405),
            .in2(N__2495),
            .in3(N__2475),
            .lcout(ctrl_tap_instruction_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4313),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_tap_instruction_i2_LC_5_5_5.C_ON=1'b0;
    defparam ctrl_tap_instruction_i2_LC_5_5_5.SEQ_MODE=4'b1000;
    defparam ctrl_tap_instruction_i2_LC_5_5_5.LUT_INIT=16'b1111011110110011;
    LogicCell40 ctrl_tap_instruction_i2_LC_5_5_5 (
            .in0(N__2404),
            .in1(N__3204),
            .in2(N__2447),
            .in3(N__2432),
            .lcout(ctrl_tap_instruction_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4313),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_tap_instruction_i1_LC_5_5_6.C_ON=1'b0;
    defparam ctrl_tap_instruction_i1_LC_5_5_6.SEQ_MODE=4'b1000;
    defparam ctrl_tap_instruction_i1_LC_5_5_6.LUT_INIT=16'b1010001010000000;
    LogicCell40 ctrl_tap_instruction_i1_LC_5_5_6 (
            .in0(N__3203),
            .in1(N__2403),
            .in2(N__2393),
            .in3(N__2376),
            .lcout(ctrl_tap_instruction_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4313),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_tap_fsm_state_i1_LC_5_5_7.C_ON=1'b0;
    defparam ctrl_tap_fsm_state_i1_LC_5_5_7.SEQ_MODE=4'b1000;
    defparam ctrl_tap_fsm_state_i1_LC_5_5_7.LUT_INIT=16'b1111100000001000;
    LogicCell40 ctrl_tap_fsm_state_i1_LC_5_5_7 (
            .in0(N__4204),
            .in1(N__2345),
            .in2(N__4235),
            .in3(N__3608),
            .lcout(ctrl_tap_fsm_state_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4313),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_1_LC_5_6_0.C_ON=1'b0;
    defparam i1_2_lut_adj_1_LC_5_6_0.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_1_LC_5_6_0.LUT_INIT=16'b1010101000000000;
    LogicCell40 i1_2_lut_adj_1_LC_5_6_0 (
            .in0(N__3821),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4120),
            .lcout(),
            .ltout(n118_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1539_2_lut_3_lut_4_lut_LC_5_6_1.C_ON=1'b0;
    defparam i1539_2_lut_3_lut_4_lut_LC_5_6_1.SEQ_MODE=4'b0000;
    defparam i1539_2_lut_3_lut_4_lut_LC_5_6_1.LUT_INIT=16'b1110111111111111;
    LogicCell40 i1539_2_lut_3_lut_4_lut_LC_5_6_1 (
            .in0(N__3707),
            .in1(N__3952),
            .in2(N__2339),
            .in3(N__4023),
            .lcout(n2273),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1531_3_lut_4_lut_LC_5_6_2.C_ON=1'b0;
    defparam i1531_3_lut_4_lut_LC_5_6_2.SEQ_MODE=4'b0000;
    defparam i1531_3_lut_4_lut_LC_5_6_2.LUT_INIT=16'b0111011101100111;
    LogicCell40 i1531_3_lut_4_lut_LC_5_6_2 (
            .in0(N__3822),
            .in1(N__3951),
            .in2(N__4042),
            .in3(N__4121),
            .lcout(),
            .ltout(n2282_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n2323_bdd_4_lut_LC_5_6_3.C_ON=1'b0;
    defparam n2323_bdd_4_lut_LC_5_6_3.SEQ_MODE=4'b0000;
    defparam n2323_bdd_4_lut_LC_5_6_3.LUT_INIT=16'b1100110010111000;
    LogicCell40 n2323_bdd_4_lut_LC_5_6_3 (
            .in0(N__3746),
            .in1(N__2540),
            .in2(N__2579),
            .in3(N__4202),
            .lcout(),
            .ltout(n2326_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_tap_fsm_state_i0_LC_5_6_4.C_ON=1'b0;
    defparam ctrl_tap_fsm_state_i0_LC_5_6_4.SEQ_MODE=4'b1000;
    defparam ctrl_tap_fsm_state_i0_LC_5_6_4.LUT_INIT=16'b1011000111110101;
    LogicCell40 ctrl_tap_fsm_state_i0_LC_5_6_4 (
            .in0(N__4226),
            .in1(N__3950),
            .in2(N__2576),
            .in3(N__2573),
            .lcout(ctrl_tap_fsm_state_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4310),
            .ce(),
            .sr(_gnd_net_));
    defparam i1482_4_lut_LC_5_6_5.C_ON=1'b0;
    defparam i1482_4_lut_LC_5_6_5.SEQ_MODE=4'b0000;
    defparam i1482_4_lut_LC_5_6_5.LUT_INIT=16'b1011101110111000;
    LogicCell40 i1482_4_lut_LC_5_6_5 (
            .in0(N__2534),
            .in1(N__4201),
            .in2(N__2567),
            .in3(N__4259),
            .lcout(),
            .ltout(n2231_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_tap_fsm_state_i2_LC_5_6_6.C_ON=1'b0;
    defparam ctrl_tap_fsm_state_i2_LC_5_6_6.SEQ_MODE=4'b1000;
    defparam ctrl_tap_fsm_state_i2_LC_5_6_6.LUT_INIT=16'b1110010010100000;
    LogicCell40 ctrl_tap_fsm_state_i2_LC_5_6_6 (
            .in0(N__4227),
            .in1(N__4203),
            .in2(N__2552),
            .in3(N__2549),
            .lcout(ctrl_tap_fsm_state_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4310),
            .ce(),
            .sr(_gnd_net_));
    defparam n2317_bdd_4_lut_4_lut_LC_5_6_7.C_ON=1'b0;
    defparam n2317_bdd_4_lut_4_lut_LC_5_6_7.SEQ_MODE=4'b0000;
    defparam n2317_bdd_4_lut_4_lut_LC_5_6_7.LUT_INIT=16'b0111110011100000;
    LogicCell40 n2317_bdd_4_lut_4_lut_LC_5_6_7 (
            .in0(N__3706),
            .in1(N__4022),
            .in2(N__4143),
            .in3(N__3820),
            .lcout(n1119),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1535_2_lut_3_lut_LC_5_7_0.C_ON=1'b0;
    defparam i1535_2_lut_3_lut_LC_5_7_0.SEQ_MODE=4'b0000;
    defparam i1535_2_lut_3_lut_LC_5_7_0.LUT_INIT=16'b0010001000000000;
    LogicCell40 i1535_2_lut_3_lut_LC_5_7_0 (
            .in0(N__4123),
            .in1(N__3943),
            .in2(_gnd_net_),
            .in3(N__3848),
            .lcout(),
            .ltout(n2263_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_tap_fsm_state_0__bdd_4_lut_4_lut_LC_5_7_1.C_ON=1'b0;
    defparam ctrl_tap_fsm_state_0__bdd_4_lut_4_lut_LC_5_7_1.SEQ_MODE=4'b0000;
    defparam ctrl_tap_fsm_state_0__bdd_4_lut_4_lut_LC_5_7_1.LUT_INIT=16'b1110011011000100;
    LogicCell40 ctrl_tap_fsm_state_0__bdd_4_lut_4_lut_LC_5_7_1 (
            .in0(N__4198),
            .in1(N__3719),
            .in2(N__2543),
            .in3(N__2726),
            .lcout(n2323),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1557_4_lut_4_lut_LC_5_7_2.C_ON=1'b0;
    defparam i1557_4_lut_4_lut_LC_5_7_2.SEQ_MODE=4'b0000;
    defparam i1557_4_lut_4_lut_LC_5_7_2.LUT_INIT=16'b1001110100010101;
    LogicCell40 i1557_4_lut_4_lut_LC_5_7_2 (
            .in0(N__4124),
            .in1(N__3944),
            .in2(N__3733),
            .in3(N__3849),
            .lcout(n2272),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_ledsArea_store_i0_i8_LC_5_7_3.C_ON=1'b0;
    defparam ctrl_ledsArea_store_i0_i8_LC_5_7_3.SEQ_MODE=4'b1000;
    defparam ctrl_ledsArea_store_i0_i8_LC_5_7_3.LUT_INIT=16'b1111010110100000;
    LogicCell40 ctrl_ledsArea_store_i0_i8_LC_5_7_3 (
            .in0(N__4393),
            .in1(_gnd_net_),
            .in2(N__2800),
            .in3(N__4642),
            .lcout(io_leds_c_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4308),
            .ce(),
            .sr(_gnd_net_));
    defparam i1041_4_lut_4_lut_LC_5_7_4.C_ON=1'b0;
    defparam i1041_4_lut_4_lut_LC_5_7_4.SEQ_MODE=4'b0000;
    defparam i1041_4_lut_4_lut_LC_5_7_4.LUT_INIT=16'b1101111101011110;
    LogicCell40 i1041_4_lut_4_lut_LC_5_7_4 (
            .in0(N__4036),
            .in1(N__3720),
            .in2(N__4144),
            .in3(N__3850),
            .lcout(n1117),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1473_4_lut_LC_5_7_6.C_ON=1'b0;
    defparam i1473_4_lut_LC_5_7_6.SEQ_MODE=4'b0000;
    defparam i1473_4_lut_LC_5_7_6.LUT_INIT=16'b1000000000000000;
    LogicCell40 i1473_4_lut_LC_5_7_6 (
            .in0(N__2776),
            .in1(N__2764),
            .in2(N__2753),
            .in3(N__2737),
            .lcout(n2222),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1558_2_lut_LC_5_7_7.C_ON=1'b0;
    defparam i1558_2_lut_LC_5_7_7.SEQ_MODE=4'b0000;
    defparam i1558_2_lut_LC_5_7_7.LUT_INIT=16'b0101010110101010;
    LogicCell40 i1558_2_lut_LC_5_7_7 (
            .in0(N__3945),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4122),
            .lcout(n2309),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1467_4_lut_LC_5_8_0.C_ON=1'b0;
    defparam i1467_4_lut_LC_5_8_0.SEQ_MODE=4'b0000;
    defparam i1467_4_lut_LC_5_8_0.LUT_INIT=16'b1000000000000000;
    LogicCell40 i1467_4_lut_LC_5_8_0 (
            .in0(N__2719),
            .in1(N__2707),
            .in2(N__2696),
            .in3(N__2680),
            .lcout(n2216),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1469_4_lut_LC_5_8_1.C_ON=1'b0;
    defparam i1469_4_lut_LC_5_8_1.SEQ_MODE=4'b0000;
    defparam i1469_4_lut_LC_5_8_1.LUT_INIT=16'b1000000000000000;
    LogicCell40 i1469_4_lut_LC_5_8_1 (
            .in0(N__2668),
            .in1(N__2656),
            .in2(N__2645),
            .in3(N__2629),
            .lcout(),
            .ltout(n2218_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1479_4_lut_LC_5_8_2.C_ON=1'b0;
    defparam i1479_4_lut_LC_5_8_2.SEQ_MODE=4'b0000;
    defparam i1479_4_lut_LC_5_8_2.LUT_INIT=16'b1000000000000000;
    LogicCell40 i1479_4_lut_LC_5_8_2 (
            .in0(N__2618),
            .in1(N__2948),
            .in2(N__2612),
            .in3(N__2609),
            .lcout(),
            .ltout(n2228_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i7_4_lut_LC_5_8_3.C_ON=1'b0;
    defparam i7_4_lut_LC_5_8_3.SEQ_MODE=4'b0000;
    defparam i7_4_lut_LC_5_8_3.LUT_INIT=16'b1111111111101111;
    LogicCell40 i7_4_lut_LC_5_8_3 (
            .in0(N__2602),
            .in1(N__3005),
            .in2(N__2591),
            .in3(N__2891),
            .lcout(n2185),
            .ltout(n2185_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1116_2_lut_LC_5_8_4.C_ON=1'b0;
    defparam i1116_2_lut_LC_5_8_4.SEQ_MODE=4'b0000;
    defparam i1116_2_lut_LC_5_8_4.LUT_INIT=16'b0101000001010000;
    LogicCell40 i1116_2_lut_LC_5_8_4 (
            .in0(N__2885),
            .in1(_gnd_net_),
            .in2(N__3122),
            .in3(_gnd_net_),
            .lcout(n1848),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i3_2_lut_LC_5_8_5.C_ON=1'b0;
    defparam i3_2_lut_LC_5_8_5.SEQ_MODE=4'b0000;
    defparam i3_2_lut_LC_5_8_5.LUT_INIT=16'b1111111111001100;
    LogicCell40 i3_2_lut_LC_5_8_5 (
            .in0(_gnd_net_),
            .in1(N__3028),
            .in2(_gnd_net_),
            .in3(N__3016),
            .lcout(n11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1471_4_lut_LC_5_9_0.C_ON=1'b0;
    defparam i1471_4_lut_LC_5_9_0.SEQ_MODE=4'b0000;
    defparam i1471_4_lut_LC_5_9_0.LUT_INIT=16'b1000000000000000;
    LogicCell40 i1471_4_lut_LC_5_9_0 (
            .in0(N__2998),
            .in1(N__2986),
            .in2(N__2975),
            .in3(N__2959),
            .lcout(n2220),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i5_4_lut_LC_5_9_4.C_ON=1'b0;
    defparam i5_4_lut_LC_5_9_4.SEQ_MODE=4'b0000;
    defparam i5_4_lut_LC_5_9_4.LUT_INIT=16'b1111111111111110;
    LogicCell40 i5_4_lut_LC_5_9_4 (
            .in0(N__2941),
            .in1(N__2929),
            .in2(N__2918),
            .in3(N__2902),
            .lcout(n13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_ledsArea_store_i0_i7_LC_5_9_6.C_ON=1'b0;
    defparam ctrl_ledsArea_store_i0_i7_LC_5_9_6.SEQ_MODE=4'b1000;
    defparam ctrl_ledsArea_store_i0_i7_LC_5_9_6.LUT_INIT=16'b1101110110001000;
    LogicCell40 ctrl_ledsArea_store_i0_i7_LC_5_9_6 (
            .in0(N__4414),
            .in1(N__4582),
            .in2(_gnd_net_),
            .in3(N__4520),
            .lcout(io_leds_c_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4304),
            .ce(),
            .sr(_gnd_net_));
    defparam myClockArea_toggle_92_LC_5_11_6.C_ON=1'b0;
    defparam myClockArea_toggle_92_LC_5_11_6.SEQ_MODE=4'b1000;
    defparam myClockArea_toggle_92_LC_5_11_6.LUT_INIT=16'b0011001111001100;
    LogicCell40 myClockArea_toggle_92_LC_5_11_6 (
            .in0(_gnd_net_),
            .in1(N__2860),
            .in2(_gnd_net_),
            .in3(N__2884),
            .lcout(io_leds_c_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2849),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_idcodeArea_shifter_i24_LC_6_3_1.C_ON=1'b0;
    defparam ctrl_idcodeArea_shifter_i24_LC_6_3_1.SEQ_MODE=4'b1000;
    defparam ctrl_idcodeArea_shifter_i24_LC_6_3_1.LUT_INIT=16'b1101111110001111;
    LogicCell40 ctrl_idcodeArea_shifter_i24_LC_6_3_1 (
            .in0(N__3428),
            .in1(N__2818),
            .in2(N__3299),
            .in3(N__2827),
            .lcout(ctrl_idcodeArea_shifter_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4321),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_idcodeArea_shifter_i25_LC_6_3_2.C_ON=1'b0;
    defparam ctrl_idcodeArea_shifter_i25_LC_6_3_2.SEQ_MODE=4'b1000;
    defparam ctrl_idcodeArea_shifter_i25_LC_6_3_2.LUT_INIT=16'b1011101111110011;
    LogicCell40 ctrl_idcodeArea_shifter_i25_LC_6_3_2 (
            .in0(N__2828),
            .in1(N__3290),
            .in2(N__3538),
            .in3(N__3429),
            .lcout(ctrl_idcodeArea_shifter_25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4321),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_idcodeArea_shifter_i23_LC_6_3_4.C_ON=1'b0;
    defparam ctrl_idcodeArea_shifter_i23_LC_6_3_4.SEQ_MODE=4'b1000;
    defparam ctrl_idcodeArea_shifter_i23_LC_6_3_4.LUT_INIT=16'b1000100011000000;
    LogicCell40 ctrl_idcodeArea_shifter_i23_LC_6_3_4 (
            .in0(N__3484),
            .in1(N__3286),
            .in2(N__2819),
            .in3(N__3427),
            .lcout(ctrl_idcodeArea_shifter_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4321),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_idcodeArea_shifter_i26_LC_6_3_6.C_ON=1'b0;
    defparam ctrl_idcodeArea_shifter_i26_LC_6_3_6.SEQ_MODE=4'b1000;
    defparam ctrl_idcodeArea_shifter_i26_LC_6_3_6.LUT_INIT=16'b1111001110111011;
    LogicCell40 ctrl_idcodeArea_shifter_i26_LC_6_3_6 (
            .in0(N__3550),
            .in1(N__3291),
            .in2(N__3539),
            .in3(N__3430),
            .lcout(ctrl_idcodeArea_shifter_26),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4321),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_tap_bypass_83_LC_6_4_0.C_ON=1'b0;
    defparam ctrl_tap_bypass_83_LC_6_4_0.SEQ_MODE=4'b1000;
    defparam ctrl_tap_bypass_83_LC_6_4_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 ctrl_tap_bypass_83_LC_6_4_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3523),
            .lcout(ctrl_tap_bypass),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4320),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_idcodeArea_shifter_i20_LC_6_4_1.C_ON=1'b0;
    defparam ctrl_idcodeArea_shifter_i20_LC_6_4_1.SEQ_MODE=4'b1000;
    defparam ctrl_idcodeArea_shifter_i20_LC_6_4_1.LUT_INIT=16'b1110010000000000;
    LogicCell40 ctrl_idcodeArea_shifter_i20_LC_6_4_1 (
            .in0(N__3411),
            .in1(N__3454),
            .in2(N__3314),
            .in3(N__3248),
            .lcout(ctrl_idcodeArea_shifter_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4320),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_idcodeArea_shifter_i22_LC_6_4_2.C_ON=1'b0;
    defparam ctrl_idcodeArea_shifter_i22_LC_6_4_2.SEQ_MODE=4'b1000;
    defparam ctrl_idcodeArea_shifter_i22_LC_6_4_2.LUT_INIT=16'b1011101111110011;
    LogicCell40 ctrl_idcodeArea_shifter_i22_LC_6_4_2 (
            .in0(N__3469),
            .in1(N__3246),
            .in2(N__3485),
            .in3(N__3413),
            .lcout(ctrl_idcodeArea_shifter_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4320),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_idcodeArea_shifter_i21_LC_6_4_3.C_ON=1'b0;
    defparam ctrl_idcodeArea_shifter_i21_LC_6_4_3.SEQ_MODE=4'b1000;
    defparam ctrl_idcodeArea_shifter_i21_LC_6_4_3.LUT_INIT=16'b1101100011111111;
    LogicCell40 ctrl_idcodeArea_shifter_i21_LC_6_4_3 (
            .in0(N__3412),
            .in1(N__3455),
            .in2(N__3470),
            .in3(N__3249),
            .lcout(ctrl_idcodeArea_shifter_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4320),
            .ce(),
            .sr(_gnd_net_));
    defparam i1017_3_lut_4_lut_LC_6_4_4.C_ON=1'b0;
    defparam i1017_3_lut_4_lut_LC_6_4_4.SEQ_MODE=4'b0000;
    defparam i1017_3_lut_4_lut_LC_6_4_4.LUT_INIT=16'b1110101001101010;
    LogicCell40 i1017_3_lut_4_lut_LC_6_4_4 (
            .in0(N__4152),
            .in1(N__3731),
            .in2(N__3949),
            .in3(N__3840),
            .lcout(n929),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_idcodeArea_shifter_i18_LC_6_4_6.C_ON=1'b0;
    defparam ctrl_idcodeArea_shifter_i18_LC_6_4_6.SEQ_MODE=4'b1000;
    defparam ctrl_idcodeArea_shifter_i18_LC_6_4_6.LUT_INIT=16'b1011101111110011;
    LogicCell40 ctrl_idcodeArea_shifter_i18_LC_6_4_6 (
            .in0(N__3445),
            .in1(N__3245),
            .in2(N__3134),
            .in3(N__3409),
            .lcout(ctrl_idcodeArea_shifter_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4320),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_idcodeArea_shifter_i19_LC_6_4_7.C_ON=1'b0;
    defparam ctrl_idcodeArea_shifter_i19_LC_6_4_7.SEQ_MODE=4'b1000;
    defparam ctrl_idcodeArea_shifter_i19_LC_6_4_7.LUT_INIT=16'b1101100000000000;
    LogicCell40 ctrl_idcodeArea_shifter_i19_LC_6_4_7 (
            .in0(N__3410),
            .in1(N__3133),
            .in2(N__3313),
            .in3(N__3247),
            .lcout(ctrl_idcodeArea_shifter_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4320),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_LC_6_5_0.C_ON=1'b0;
    defparam i1_2_lut_LC_6_5_0.SEQ_MODE=4'b0000;
    defparam i1_2_lut_LC_6_5_0.LUT_INIT=16'b0011001100000000;
    LogicCell40 i1_2_lut_LC_6_5_0 (
            .in0(_gnd_net_),
            .in1(N__4110),
            .in2(_gnd_net_),
            .in3(N__4017),
            .lcout(n4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_adj_4_LC_6_5_1.C_ON=1'b0;
    defparam i1_2_lut_3_lut_adj_4_LC_6_5_1.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_adj_4_LC_6_5_1.LUT_INIT=16'b1111111111111010;
    LogicCell40 i1_2_lut_3_lut_adj_4_LC_6_5_1 (
            .in0(N__4021),
            .in1(_gnd_net_),
            .in2(N__3955),
            .in3(N__4153),
            .lcout(),
            .ltout(n17_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i954_4_lut_LC_6_5_2.C_ON=1'b0;
    defparam i954_4_lut_LC_6_5_2.SEQ_MODE=4'b0000;
    defparam i954_4_lut_LC_6_5_2.LUT_INIT=16'b1100110000001010;
    LogicCell40 i954_4_lut_LC_6_5_2 (
            .in0(N__3817),
            .in1(N__4258),
            .in2(N__3614),
            .in3(N__3698),
            .lcout(),
            .ltout(n1687_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1485_3_lut_LC_6_5_3.C_ON=1'b0;
    defparam i1485_3_lut_LC_6_5_3.SEQ_MODE=4'b0000;
    defparam i1485_3_lut_LC_6_5_3.LUT_INIT=16'b0011001111110000;
    LogicCell40 i1485_3_lut_LC_6_5_3 (
            .in0(_gnd_net_),
            .in1(N__3602),
            .in2(N__3611),
            .in3(N__4200),
            .lcout(n2234),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i13_4_lut_LC_6_5_4.C_ON=1'b0;
    defparam i13_4_lut_LC_6_5_4.SEQ_MODE=4'b0000;
    defparam i13_4_lut_LC_6_5_4.LUT_INIT=16'b1000100011110000;
    LogicCell40 i13_4_lut_LC_6_5_4 (
            .in0(N__3816),
            .in1(N__3939),
            .in2(N__3730),
            .in3(N__4112),
            .lcout(n8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_3_lut_4_lut_LC_6_5_5.C_ON=1'b0;
    defparam i2_3_lut_4_lut_LC_6_5_5.SEQ_MODE=4'b0000;
    defparam i2_3_lut_4_lut_LC_6_5_5.LUT_INIT=16'b1111011111111111;
    LogicCell40 i2_3_lut_4_lut_LC_6_5_5 (
            .in0(N__4111),
            .in1(N__3815),
            .in2(N__4041),
            .in3(N__3699),
            .lcout(n7_adj_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1449_2_lut_LC_6_5_6.C_ON=1'b0;
    defparam i1449_2_lut_LC_6_5_6.SEQ_MODE=4'b0000;
    defparam i1449_2_lut_LC_6_5_6.LUT_INIT=16'b1111111110101010;
    LogicCell40 i1449_2_lut_LC_6_5_6 (
            .in0(N__3814),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3697),
            .lcout(n2198),
            .ltout(n2198_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1182_4_lut_LC_6_5_7.C_ON=1'b0;
    defparam i1182_4_lut_LC_6_5_7.SEQ_MODE=4'b0000;
    defparam i1182_4_lut_LC_6_5_7.LUT_INIT=16'b1100101011001100;
    LogicCell40 i1182_4_lut_LC_6_5_7 (
            .in0(N__3590),
            .in1(N__3575),
            .in2(N__3569),
            .in3(N__3566),
            .lcout(ctrl_tap_tdoUnbufferd_N_213),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_4_lut_adj_6_LC_6_6_0.C_ON=1'b0;
    defparam i1_2_lut_3_lut_4_lut_adj_6_LC_6_6_0.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_4_lut_adj_6_LC_6_6_0.LUT_INIT=16'b0000001000000000;
    LogicCell40 i1_2_lut_3_lut_4_lut_adj_6_LC_6_6_0 (
            .in0(N__3841),
            .in1(N__3725),
            .in2(N__4043),
            .in3(N__4115),
            .lcout(n1638),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_LC_6_6_1.C_ON=1'b0;
    defparam i1_2_lut_3_lut_LC_6_6_1.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_LC_6_6_1.LUT_INIT=16'b0010001000000000;
    LogicCell40 i1_2_lut_3_lut_LC_6_6_1 (
            .in0(N__4114),
            .in1(N__4028),
            .in2(_gnd_net_),
            .in3(N__3842),
            .lcout(n2186),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_ledsArea_store_i0_i4_LC_6_6_2.C_ON=1'b0;
    defparam ctrl_ledsArea_store_i0_i4_LC_6_6_2.SEQ_MODE=4'b1000;
    defparam ctrl_ledsArea_store_i0_i4_LC_6_6_2.LUT_INIT=16'b1010101011001100;
    LogicCell40 ctrl_ledsArea_store_i0_i4_LC_6_6_2 (
            .in0(N__4720),
            .in1(N__4709),
            .in2(_gnd_net_),
            .in3(N__4401),
            .lcout(ctrl_ledsArea_store_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4314),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_4_lut_adj_7_LC_6_6_3.C_ON=1'b0;
    defparam i1_2_lut_4_lut_adj_7_LC_6_6_3.SEQ_MODE=4'b0000;
    defparam i1_2_lut_4_lut_adj_7_LC_6_6_3.LUT_INIT=16'b0000000000000100;
    LogicCell40 i1_2_lut_4_lut_adj_7_LC_6_6_3 (
            .in0(N__4113),
            .in1(N__4027),
            .in2(N__3851),
            .in3(N__3954),
            .lcout(n1686),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_ledsArea_store_i0_i2_LC_6_6_4.C_ON=1'b0;
    defparam ctrl_ledsArea_store_i0_i2_LC_6_6_4.SEQ_MODE=4'b1000;
    defparam ctrl_ledsArea_store_i0_i2_LC_6_6_4.LUT_INIT=16'b1010101011001100;
    LogicCell40 ctrl_ledsArea_store_i0_i2_LC_6_6_4 (
            .in0(N__4755),
            .in1(N__4738),
            .in2(_gnd_net_),
            .in3(N__4400),
            .lcout(io_leds_c_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4314),
            .ce(),
            .sr(_gnd_net_));
    defparam i114_3_lut_LC_6_6_5.C_ON=1'b0;
    defparam i114_3_lut_LC_6_6_5.SEQ_MODE=4'b0000;
    defparam i114_3_lut_LC_6_6_5.LUT_INIT=16'b1100110010111011;
    LogicCell40 i114_3_lut_LC_6_6_5 (
            .in0(N__3726),
            .in1(N__4032),
            .in2(_gnd_net_),
            .in3(N__3843),
            .lcout(),
            .ltout(n112_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1534_3_lut_LC_6_6_6.C_ON=1'b0;
    defparam i1534_3_lut_LC_6_6_6.SEQ_MODE=4'b0000;
    defparam i1534_3_lut_LC_6_6_6.LUT_INIT=16'b1010101010100000;
    LogicCell40 i1534_3_lut_LC_6_6_6 (
            .in0(N__3953),
            .in1(_gnd_net_),
            .in2(N__4247),
            .in3(N__4116),
            .lcout(),
            .ltout(n2260_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_tap_fsm_state_i3_LC_6_6_7.C_ON=1'b0;
    defparam ctrl_tap_fsm_state_i3_LC_6_6_7.SEQ_MODE=4'b1000;
    defparam ctrl_tap_fsm_state_i3_LC_6_6_7.LUT_INIT=16'b1011101111000000;
    LogicCell40 ctrl_tap_fsm_state_i3_LC_6_6_7 (
            .in0(N__4244),
            .in1(N__4231),
            .in2(N__4208),
            .in3(N__4205),
            .lcout(ctrl_tap_fsm_state_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4314),
            .ce(),
            .sr(_gnd_net_));
    defparam i1494_3_lut_4_lut_LC_6_7_4.C_ON=1'b0;
    defparam i1494_3_lut_4_lut_LC_6_7_4.SEQ_MODE=4'b0000;
    defparam i1494_3_lut_4_lut_LC_6_7_4.LUT_INIT=16'b1111111010111011;
    LogicCell40 i1494_3_lut_4_lut_LC_6_7_4 (
            .in0(N__4142),
            .in1(N__4037),
            .in2(N__3956),
            .in3(N__3847),
            .lcout(n2243),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_ledsArea_shifter_i0_i4_LC_7_6_0.C_ON=1'b0;
    defparam ctrl_ledsArea_shifter_i0_i4_LC_7_6_0.SEQ_MODE=4'b1000;
    defparam ctrl_ledsArea_shifter_i0_i4_LC_7_6_0.LUT_INIT=16'b1100000010001000;
    LogicCell40 ctrl_ledsArea_shifter_i0_i4_LC_7_6_0 (
            .in0(N__4450),
            .in1(N__3740),
            .in2(N__4663),
            .in3(N__3734),
            .lcout(ctrl_ledsArea_shifter_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4318),
            .ce(N__4502),
            .sr(_gnd_net_));
    defparam ctrl_ledsArea_shifter_i0_i1_LC_7_6_1.C_ON=1'b0;
    defparam ctrl_ledsArea_shifter_i0_i1_LC_7_6_1.SEQ_MODE=4'b1000;
    defparam ctrl_ledsArea_shifter_i0_i1_LC_7_6_1.LUT_INIT=16'b1100000010101010;
    LogicCell40 ctrl_ledsArea_shifter_i0_i1_LC_7_6_1 (
            .in0(N__4429),
            .in1(N__4624),
            .in2(N__4762),
            .in3(N__4553),
            .lcout(ctrl_ledsArea_shifter_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4318),
            .ce(N__4502),
            .sr(_gnd_net_));
    defparam ctrl_ledsArea_shifter_i0_i2_LC_7_6_2.C_ON=1'b0;
    defparam ctrl_ledsArea_shifter_i0_i2_LC_7_6_2.SEQ_MODE=4'b1000;
    defparam ctrl_ledsArea_shifter_i0_i2_LC_7_6_2.LUT_INIT=16'b1110010001000100;
    LogicCell40 ctrl_ledsArea_shifter_i0_i2_LC_7_6_2 (
            .in0(N__4554),
            .in1(N__4708),
            .in2(N__4351),
            .in3(N__4627),
            .lcout(ctrl_ledsArea_shifter_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4318),
            .ce(N__4502),
            .sr(_gnd_net_));
    defparam ctrl_ledsArea_shifter_i0_i3_LC_7_6_3.C_ON=1'b0;
    defparam ctrl_ledsArea_shifter_i0_i3_LC_7_6_3.SEQ_MODE=4'b1000;
    defparam ctrl_ledsArea_shifter_i0_i3_LC_7_6_3.LUT_INIT=16'b1100000010101010;
    LogicCell40 ctrl_ledsArea_shifter_i0_i3_LC_7_6_3 (
            .in0(N__4472),
            .in1(N__4625),
            .in2(N__4724),
            .in3(N__4555),
            .lcout(ctrl_ledsArea_shifter_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4318),
            .ce(N__4502),
            .sr(_gnd_net_));
    defparam ctrl_ledsArea_shifter_i0_i5_LC_7_6_4.C_ON=1'b0;
    defparam ctrl_ledsArea_shifter_i0_i5_LC_7_6_4.SEQ_MODE=4'b1000;
    defparam ctrl_ledsArea_shifter_i0_i5_LC_7_6_4.LUT_INIT=16'b1110010001000100;
    LogicCell40 ctrl_ledsArea_shifter_i0_i5_LC_7_6_4 (
            .in0(N__4556),
            .in1(N__4513),
            .in2(N__4696),
            .in3(N__4628),
            .lcout(ctrl_ledsArea_shifter_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4318),
            .ce(N__4502),
            .sr(_gnd_net_));
    defparam ctrl_ledsArea_shifter_i0_i6_LC_7_6_5.C_ON=1'b0;
    defparam ctrl_ledsArea_shifter_i0_i6_LC_7_6_5.SEQ_MODE=4'b1000;
    defparam ctrl_ledsArea_shifter_i0_i6_LC_7_6_5.LUT_INIT=16'b1100000010101010;
    LogicCell40 ctrl_ledsArea_shifter_i0_i6_LC_7_6_5 (
            .in0(N__4643),
            .in1(N__4626),
            .in2(N__4600),
            .in3(N__4557),
            .lcout(ctrl_ledsArea_shifter_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4318),
            .ce(N__4502),
            .sr(_gnd_net_));
    defparam ctrl_ledsArea_store_i0_i5_LC_7_7_2.C_ON=1'b0;
    defparam ctrl_ledsArea_store_i0_i5_LC_7_7_2.SEQ_MODE=4'b1000;
    defparam ctrl_ledsArea_store_i0_i5_LC_7_7_2.LUT_INIT=16'b1010101011001100;
    LogicCell40 ctrl_ledsArea_store_i0_i5_LC_7_7_2 (
            .in0(N__4449),
            .in1(N__4471),
            .in2(_gnd_net_),
            .in3(N__4416),
            .lcout(io_leds_c_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4315),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_ledsArea_store_i0_i3_LC_7_8_1.C_ON=1'b0;
    defparam ctrl_ledsArea_store_i0_i3_LC_7_8_1.SEQ_MODE=4'b1000;
    defparam ctrl_ledsArea_store_i0_i3_LC_7_8_1.LUT_INIT=16'b1010101011001100;
    LogicCell40 ctrl_ledsArea_store_i0_i3_LC_7_8_1 (
            .in0(N__4338),
            .in1(N__4433),
            .in2(_gnd_net_),
            .in3(N__4417),
            .lcout(io_leds_c_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4311),
            .ce(),
            .sr(_gnd_net_));
endmodule // MyTopLevel
