// ******************************************************************************

// iCEcube Netlister

// Version:            2017.08.27940

// Build Date:         Sep 12 2017 08:25:46

// File Generated:     Apr 28 2020 10:13:15

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "MyTopLevel" view "INTERFACE"

module MyTopLevel (
    io_leds,
    io_jtag_tms,
    io_jtag_tdo,
    io_jtag_tdi,
    io_jtag_tck,
    global_reset,
    global_clk);

    output [7:0] io_leds;
    input io_jtag_tms;
    output io_jtag_tdo;
    input io_jtag_tdi;
    input io_jtag_tck;
    input global_reset;
    input global_clk;

    wire N__5400;
    wire N__5399;
    wire N__5398;
    wire N__5389;
    wire N__5388;
    wire N__5387;
    wire N__5380;
    wire N__5379;
    wire N__5378;
    wire N__5371;
    wire N__5370;
    wire N__5369;
    wire N__5362;
    wire N__5361;
    wire N__5360;
    wire N__5353;
    wire N__5352;
    wire N__5351;
    wire N__5344;
    wire N__5343;
    wire N__5342;
    wire N__5335;
    wire N__5334;
    wire N__5333;
    wire N__5326;
    wire N__5325;
    wire N__5324;
    wire N__5317;
    wire N__5316;
    wire N__5315;
    wire N__5308;
    wire N__5307;
    wire N__5306;
    wire N__5299;
    wire N__5298;
    wire N__5297;
    wire N__5290;
    wire N__5289;
    wire N__5288;
    wire N__5281;
    wire N__5280;
    wire N__5279;
    wire N__5262;
    wire N__5261;
    wire N__5258;
    wire N__5257;
    wire N__5254;
    wire N__5251;
    wire N__5248;
    wire N__5245;
    wire N__5238;
    wire N__5235;
    wire N__5232;
    wire N__5229;
    wire N__5228;
    wire N__5225;
    wire N__5222;
    wire N__5217;
    wire N__5216;
    wire N__5215;
    wire N__5214;
    wire N__5213;
    wire N__5202;
    wire N__5199;
    wire N__5196;
    wire N__5195;
    wire N__5192;
    wire N__5189;
    wire N__5186;
    wire N__5185;
    wire N__5182;
    wire N__5181;
    wire N__5178;
    wire N__5175;
    wire N__5172;
    wire N__5169;
    wire N__5164;
    wire N__5157;
    wire N__5154;
    wire N__5151;
    wire N__5148;
    wire N__5145;
    wire N__5144;
    wire N__5141;
    wire N__5138;
    wire N__5133;
    wire N__5132;
    wire N__5127;
    wire N__5124;
    wire N__5121;
    wire N__5120;
    wire N__5115;
    wire N__5112;
    wire N__5109;
    wire N__5106;
    wire N__5103;
    wire N__5102;
    wire N__5099;
    wire N__5096;
    wire N__5091;
    wire N__5090;
    wire N__5085;
    wire N__5082;
    wire N__5079;
    wire N__5078;
    wire N__5077;
    wire N__5076;
    wire N__5075;
    wire N__5074;
    wire N__5071;
    wire N__5068;
    wire N__5065;
    wire N__5064;
    wire N__5063;
    wire N__5062;
    wire N__5061;
    wire N__5058;
    wire N__5057;
    wire N__5056;
    wire N__5055;
    wire N__5054;
    wire N__5053;
    wire N__5052;
    wire N__5051;
    wire N__5050;
    wire N__5049;
    wire N__5048;
    wire N__5047;
    wire N__5046;
    wire N__5045;
    wire N__5044;
    wire N__5043;
    wire N__5042;
    wire N__5041;
    wire N__5040;
    wire N__5039;
    wire N__5038;
    wire N__5037;
    wire N__5032;
    wire N__5027;
    wire N__5024;
    wire N__5021;
    wire N__5014;
    wire N__5011;
    wire N__5002;
    wire N__4991;
    wire N__4986;
    wire N__4979;
    wire N__4968;
    wire N__4963;
    wire N__4956;
    wire N__4951;
    wire N__4944;
    wire N__4929;
    wire N__4928;
    wire N__4927;
    wire N__4926;
    wire N__4925;
    wire N__4924;
    wire N__4923;
    wire N__4922;
    wire N__4921;
    wire N__4920;
    wire N__4919;
    wire N__4918;
    wire N__4917;
    wire N__4916;
    wire N__4915;
    wire N__4914;
    wire N__4913;
    wire N__4912;
    wire N__4911;
    wire N__4910;
    wire N__4907;
    wire N__4906;
    wire N__4905;
    wire N__4904;
    wire N__4901;
    wire N__4900;
    wire N__4899;
    wire N__4898;
    wire N__4897;
    wire N__4896;
    wire N__4885;
    wire N__4878;
    wire N__4877;
    wire N__4874;
    wire N__4871;
    wire N__4870;
    wire N__4867;
    wire N__4866;
    wire N__4865;
    wire N__4864;
    wire N__4863;
    wire N__4860;
    wire N__4859;
    wire N__4858;
    wire N__4857;
    wire N__4856;
    wire N__4855;
    wire N__4854;
    wire N__4851;
    wire N__4848;
    wire N__4841;
    wire N__4832;
    wire N__4825;
    wire N__4822;
    wire N__4815;
    wire N__4810;
    wire N__4807;
    wire N__4804;
    wire N__4801;
    wire N__4796;
    wire N__4791;
    wire N__4786;
    wire N__4779;
    wire N__4770;
    wire N__4767;
    wire N__4758;
    wire N__4751;
    wire N__4728;
    wire N__4727;
    wire N__4724;
    wire N__4719;
    wire N__4716;
    wire N__4715;
    wire N__4714;
    wire N__4713;
    wire N__4712;
    wire N__4711;
    wire N__4710;
    wire N__4709;
    wire N__4708;
    wire N__4707;
    wire N__4706;
    wire N__4705;
    wire N__4704;
    wire N__4703;
    wire N__4702;
    wire N__4701;
    wire N__4700;
    wire N__4665;
    wire N__4662;
    wire N__4659;
    wire N__4656;
    wire N__4653;
    wire N__4650;
    wire N__4649;
    wire N__4646;
    wire N__4643;
    wire N__4640;
    wire N__4637;
    wire N__4636;
    wire N__4631;
    wire N__4628;
    wire N__4623;
    wire N__4622;
    wire N__4619;
    wire N__4616;
    wire N__4613;
    wire N__4610;
    wire N__4605;
    wire N__4602;
    wire N__4599;
    wire N__4596;
    wire N__4595;
    wire N__4592;
    wire N__4589;
    wire N__4588;
    wire N__4583;
    wire N__4580;
    wire N__4575;
    wire N__4572;
    wire N__4571;
    wire N__4568;
    wire N__4565;
    wire N__4560;
    wire N__4557;
    wire N__4554;
    wire N__4551;
    wire N__4548;
    wire N__4545;
    wire N__4544;
    wire N__4541;
    wire N__4538;
    wire N__4537;
    wire N__4532;
    wire N__4529;
    wire N__4524;
    wire N__4521;
    wire N__4520;
    wire N__4517;
    wire N__4514;
    wire N__4511;
    wire N__4508;
    wire N__4503;
    wire N__4500;
    wire N__4497;
    wire N__4496;
    wire N__4493;
    wire N__4490;
    wire N__4485;
    wire N__4482;
    wire N__4481;
    wire N__4478;
    wire N__4475;
    wire N__4472;
    wire N__4469;
    wire N__4464;
    wire N__4461;
    wire N__4458;
    wire N__4457;
    wire N__4454;
    wire N__4451;
    wire N__4450;
    wire N__4447;
    wire N__4444;
    wire N__4441;
    wire N__4434;
    wire N__4431;
    wire N__4428;
    wire N__4427;
    wire N__4424;
    wire N__4421;
    wire N__4416;
    wire N__4413;
    wire N__4412;
    wire N__4409;
    wire N__4408;
    wire N__4405;
    wire N__4402;
    wire N__4399;
    wire N__4392;
    wire N__4389;
    wire N__4388;
    wire N__4385;
    wire N__4382;
    wire N__4379;
    wire N__4376;
    wire N__4371;
    wire N__4368;
    wire N__4367;
    wire N__4366;
    wire N__4365;
    wire N__4364;
    wire N__4363;
    wire N__4362;
    wire N__4361;
    wire N__4358;
    wire N__4343;
    wire N__4342;
    wire N__4341;
    wire N__4338;
    wire N__4335;
    wire N__4330;
    wire N__4323;
    wire N__4320;
    wire N__4317;
    wire N__4314;
    wire N__4313;
    wire N__4310;
    wire N__4307;
    wire N__4306;
    wire N__4303;
    wire N__4300;
    wire N__4297;
    wire N__4290;
    wire N__4289;
    wire N__4288;
    wire N__4287;
    wire N__4286;
    wire N__4285;
    wire N__4284;
    wire N__4283;
    wire N__4274;
    wire N__4265;
    wire N__4260;
    wire N__4257;
    wire N__4254;
    wire N__4253;
    wire N__4250;
    wire N__4247;
    wire N__4244;
    wire N__4241;
    wire N__4236;
    wire N__4233;
    wire N__4230;
    wire N__4227;
    wire N__4224;
    wire N__4223;
    wire N__4222;
    wire N__4221;
    wire N__4220;
    wire N__4219;
    wire N__4218;
    wire N__4217;
    wire N__4216;
    wire N__4215;
    wire N__4214;
    wire N__4213;
    wire N__4210;
    wire N__4195;
    wire N__4192;
    wire N__4189;
    wire N__4188;
    wire N__4185;
    wire N__4184;
    wire N__4183;
    wire N__4182;
    wire N__4179;
    wire N__4178;
    wire N__4177;
    wire N__4176;
    wire N__4175;
    wire N__4174;
    wire N__4173;
    wire N__4172;
    wire N__4171;
    wire N__4170;
    wire N__4169;
    wire N__4168;
    wire N__4161;
    wire N__4158;
    wire N__4151;
    wire N__4148;
    wire N__4147;
    wire N__4146;
    wire N__4141;
    wire N__4138;
    wire N__4127;
    wire N__4116;
    wire N__4111;
    wire N__4106;
    wire N__4101;
    wire N__4086;
    wire N__4085;
    wire N__4084;
    wire N__4083;
    wire N__4080;
    wire N__4077;
    wire N__4076;
    wire N__4073;
    wire N__4072;
    wire N__4071;
    wire N__4070;
    wire N__4069;
    wire N__4068;
    wire N__4067;
    wire N__4066;
    wire N__4065;
    wire N__4064;
    wire N__4063;
    wire N__4062;
    wire N__4059;
    wire N__4054;
    wire N__4053;
    wire N__4052;
    wire N__4051;
    wire N__4048;
    wire N__4045;
    wire N__4042;
    wire N__4039;
    wire N__4038;
    wire N__4033;
    wire N__4030;
    wire N__4023;
    wire N__4014;
    wire N__4011;
    wire N__4004;
    wire N__3997;
    wire N__3992;
    wire N__3975;
    wire N__3974;
    wire N__3973;
    wire N__3972;
    wire N__3969;
    wire N__3968;
    wire N__3965;
    wire N__3964;
    wire N__3963;
    wire N__3962;
    wire N__3961;
    wire N__3958;
    wire N__3955;
    wire N__3950;
    wire N__3945;
    wire N__3938;
    wire N__3937;
    wire N__3934;
    wire N__3933;
    wire N__3930;
    wire N__3923;
    wire N__3920;
    wire N__3917;
    wire N__3914;
    wire N__3909;
    wire N__3906;
    wire N__3903;
    wire N__3900;
    wire N__3897;
    wire N__3894;
    wire N__3889;
    wire N__3882;
    wire N__3881;
    wire N__3880;
    wire N__3875;
    wire N__3872;
    wire N__3871;
    wire N__3870;
    wire N__3869;
    wire N__3868;
    wire N__3865;
    wire N__3864;
    wire N__3863;
    wire N__3862;
    wire N__3861;
    wire N__3860;
    wire N__3859;
    wire N__3858;
    wire N__3857;
    wire N__3856;
    wire N__3855;
    wire N__3854;
    wire N__3853;
    wire N__3850;
    wire N__3843;
    wire N__3840;
    wire N__3839;
    wire N__3838;
    wire N__3835;
    wire N__3832;
    wire N__3829;
    wire N__3818;
    wire N__3807;
    wire N__3800;
    wire N__3795;
    wire N__3780;
    wire N__3777;
    wire N__3774;
    wire N__3771;
    wire N__3768;
    wire N__3765;
    wire N__3762;
    wire N__3761;
    wire N__3758;
    wire N__3755;
    wire N__3750;
    wire N__3747;
    wire N__3746;
    wire N__3741;
    wire N__3738;
    wire N__3737;
    wire N__3734;
    wire N__3729;
    wire N__3726;
    wire N__3725;
    wire N__3720;
    wire N__3717;
    wire N__3716;
    wire N__3713;
    wire N__3710;
    wire N__3707;
    wire N__3702;
    wire N__3701;
    wire N__3698;
    wire N__3695;
    wire N__3694;
    wire N__3693;
    wire N__3692;
    wire N__3691;
    wire N__3690;
    wire N__3685;
    wire N__3684;
    wire N__3683;
    wire N__3682;
    wire N__3681;
    wire N__3678;
    wire N__3677;
    wire N__3674;
    wire N__3671;
    wire N__3670;
    wire N__3667;
    wire N__3664;
    wire N__3663;
    wire N__3660;
    wire N__3659;
    wire N__3658;
    wire N__3653;
    wire N__3650;
    wire N__3649;
    wire N__3646;
    wire N__3641;
    wire N__3636;
    wire N__3627;
    wire N__3624;
    wire N__3619;
    wire N__3614;
    wire N__3609;
    wire N__3594;
    wire N__3591;
    wire N__3590;
    wire N__3587;
    wire N__3584;
    wire N__3579;
    wire N__3576;
    wire N__3573;
    wire N__3570;
    wire N__3567;
    wire N__3566;
    wire N__3563;
    wire N__3560;
    wire N__3555;
    wire N__3554;
    wire N__3549;
    wire N__3546;
    wire N__3543;
    wire N__3540;
    wire N__3539;
    wire N__3536;
    wire N__3533;
    wire N__3532;
    wire N__3529;
    wire N__3526;
    wire N__3523;
    wire N__3520;
    wire N__3515;
    wire N__3510;
    wire N__3509;
    wire N__3506;
    wire N__3503;
    wire N__3500;
    wire N__3497;
    wire N__3494;
    wire N__3491;
    wire N__3486;
    wire N__3485;
    wire N__3482;
    wire N__3479;
    wire N__3478;
    wire N__3475;
    wire N__3472;
    wire N__3469;
    wire N__3464;
    wire N__3463;
    wire N__3460;
    wire N__3457;
    wire N__3454;
    wire N__3451;
    wire N__3448;
    wire N__3445;
    wire N__3442;
    wire N__3435;
    wire N__3432;
    wire N__3431;
    wire N__3430;
    wire N__3429;
    wire N__3428;
    wire N__3425;
    wire N__3422;
    wire N__3417;
    wire N__3414;
    wire N__3405;
    wire N__3404;
    wire N__3401;
    wire N__3398;
    wire N__3397;
    wire N__3396;
    wire N__3393;
    wire N__3390;
    wire N__3387;
    wire N__3384;
    wire N__3375;
    wire N__3372;
    wire N__3371;
    wire N__3368;
    wire N__3365;
    wire N__3360;
    wire N__3359;
    wire N__3356;
    wire N__3353;
    wire N__3352;
    wire N__3347;
    wire N__3344;
    wire N__3339;
    wire N__3336;
    wire N__3335;
    wire N__3334;
    wire N__3331;
    wire N__3326;
    wire N__3321;
    wire N__3318;
    wire N__3315;
    wire N__3312;
    wire N__3311;
    wire N__3308;
    wire N__3305;
    wire N__3300;
    wire N__3299;
    wire N__3296;
    wire N__3293;
    wire N__3292;
    wire N__3291;
    wire N__3288;
    wire N__3285;
    wire N__3280;
    wire N__3273;
    wire N__3270;
    wire N__3267;
    wire N__3264;
    wire N__3263;
    wire N__3260;
    wire N__3257;
    wire N__3252;
    wire N__3251;
    wire N__3248;
    wire N__3247;
    wire N__3244;
    wire N__3243;
    wire N__3240;
    wire N__3237;
    wire N__3232;
    wire N__3225;
    wire N__3222;
    wire N__3219;
    wire N__3218;
    wire N__3215;
    wire N__3212;
    wire N__3207;
    wire N__3204;
    wire N__3203;
    wire N__3200;
    wire N__3197;
    wire N__3192;
    wire N__3189;
    wire N__3188;
    wire N__3187;
    wire N__3186;
    wire N__3183;
    wire N__3176;
    wire N__3171;
    wire N__3168;
    wire N__3165;
    wire N__3164;
    wire N__3161;
    wire N__3158;
    wire N__3153;
    wire N__3150;
    wire N__3147;
    wire N__3146;
    wire N__3143;
    wire N__3140;
    wire N__3135;
    wire N__3132;
    wire N__3129;
    wire N__3128;
    wire N__3127;
    wire N__3126;
    wire N__3125;
    wire N__3122;
    wire N__3119;
    wire N__3116;
    wire N__3113;
    wire N__3110;
    wire N__3099;
    wire N__3096;
    wire N__3093;
    wire N__3092;
    wire N__3089;
    wire N__3086;
    wire N__3081;
    wire N__3078;
    wire N__3075;
    wire N__3074;
    wire N__3069;
    wire N__3066;
    wire N__3065;
    wire N__3060;
    wire N__3057;
    wire N__3056;
    wire N__3053;
    wire N__3050;
    wire N__3045;
    wire N__3044;
    wire N__3041;
    wire N__3038;
    wire N__3033;
    wire N__3032;
    wire N__3029;
    wire N__3026;
    wire N__3023;
    wire N__3018;
    wire N__3017;
    wire N__3014;
    wire N__3011;
    wire N__3006;
    wire N__3005;
    wire N__3002;
    wire N__2999;
    wire N__2994;
    wire N__2993;
    wire N__2990;
    wire N__2987;
    wire N__2982;
    wire N__2981;
    wire N__2978;
    wire N__2975;
    wire N__2972;
    wire N__2967;
    wire N__2966;
    wire N__2963;
    wire N__2960;
    wire N__2955;
    wire N__2952;
    wire N__2949;
    wire N__2946;
    wire N__2943;
    wire N__2940;
    wire N__2939;
    wire N__2936;
    wire N__2933;
    wire N__2928;
    wire N__2925;
    wire N__2922;
    wire N__2919;
    wire N__2916;
    wire N__2913;
    wire N__2910;
    wire N__2909;
    wire N__2908;
    wire N__2907;
    wire N__2906;
    wire N__2905;
    wire N__2904;
    wire N__2903;
    wire N__2902;
    wire N__2901;
    wire N__2900;
    wire N__2899;
    wire N__2890;
    wire N__2881;
    wire N__2880;
    wire N__2879;
    wire N__2878;
    wire N__2877;
    wire N__2876;
    wire N__2875;
    wire N__2874;
    wire N__2873;
    wire N__2872;
    wire N__2871;
    wire N__2870;
    wire N__2861;
    wire N__2858;
    wire N__2855;
    wire N__2846;
    wire N__2839;
    wire N__2830;
    wire N__2817;
    wire N__2816;
    wire N__2813;
    wire N__2810;
    wire N__2805;
    wire N__2804;
    wire N__2801;
    wire N__2798;
    wire N__2793;
    wire N__2792;
    wire N__2789;
    wire N__2786;
    wire N__2783;
    wire N__2778;
    wire N__2777;
    wire N__2774;
    wire N__2771;
    wire N__2766;
    wire N__2763;
    wire N__2760;
    wire N__2757;
    wire N__2754;
    wire N__2753;
    wire N__2752;
    wire N__2751;
    wire N__2750;
    wire N__2749;
    wire N__2748;
    wire N__2737;
    wire N__2734;
    wire N__2731;
    wire N__2724;
    wire N__2723;
    wire N__2722;
    wire N__2721;
    wire N__2712;
    wire N__2709;
    wire N__2706;
    wire N__2703;
    wire N__2702;
    wire N__2699;
    wire N__2696;
    wire N__2691;
    wire N__2690;
    wire N__2687;
    wire N__2684;
    wire N__2679;
    wire N__2678;
    wire N__2675;
    wire N__2672;
    wire N__2669;
    wire N__2664;
    wire N__2663;
    wire N__2660;
    wire N__2657;
    wire N__2652;
    wire N__2651;
    wire N__2648;
    wire N__2645;
    wire N__2640;
    wire N__2639;
    wire N__2636;
    wire N__2633;
    wire N__2630;
    wire N__2625;
    wire N__2624;
    wire N__2621;
    wire N__2618;
    wire N__2615;
    wire N__2610;
    wire N__2609;
    wire N__2606;
    wire N__2603;
    wire N__2598;
    wire N__2597;
    wire N__2594;
    wire N__2591;
    wire N__2588;
    wire N__2583;
    wire N__2582;
    wire N__2579;
    wire N__2576;
    wire N__2571;
    wire N__2570;
    wire N__2567;
    wire N__2564;
    wire N__2561;
    wire N__2556;
    wire N__2555;
    wire N__2552;
    wire N__2549;
    wire N__2546;
    wire N__2541;
    wire N__2540;
    wire N__2537;
    wire N__2532;
    wire N__2529;
    wire N__2528;
    wire N__2525;
    wire N__2522;
    wire N__2519;
    wire N__2514;
    wire N__2513;
    wire N__2512;
    wire N__2511;
    wire N__2510;
    wire N__2509;
    wire N__2508;
    wire N__2497;
    wire N__2492;
    wire N__2487;
    wire N__2486;
    wire N__2483;
    wire N__2480;
    wire N__2477;
    wire N__2472;
    wire N__2469;
    wire N__2466;
    wire N__2463;
    wire N__2460;
    wire N__2457;
    wire N__2456;
    wire N__2453;
    wire N__2450;
    wire N__2445;
    wire N__2442;
    wire N__2439;
    wire N__2438;
    wire N__2435;
    wire N__2432;
    wire N__2427;
    wire N__2424;
    wire N__2423;
    wire N__2420;
    wire N__2417;
    wire N__2412;
    wire N__2411;
    wire N__2406;
    wire N__2403;
    wire N__2400;
    wire N__2399;
    wire N__2394;
    wire N__2391;
    wire N__2388;
    wire N__2385;
    wire N__2382;
    wire N__2381;
    wire N__2378;
    wire N__2375;
    wire N__2372;
    wire N__2369;
    wire N__2364;
    wire N__2363;
    wire N__2360;
    wire N__2357;
    wire N__2354;
    wire N__2349;
    wire N__2348;
    wire N__2345;
    wire N__2342;
    wire N__2339;
    wire N__2334;
    wire N__2331;
    wire N__2330;
    wire N__2325;
    wire N__2322;
    wire N__2319;
    wire N__2318;
    wire N__2313;
    wire N__2310;
    wire N__2307;
    wire N__2306;
    wire N__2301;
    wire N__2298;
    wire N__2295;
    wire N__2292;
    wire N__2289;
    wire N__2286;
    wire N__2283;
    wire N__2280;
    wire N__2277;
    wire N__2274;
    wire N__2271;
    wire N__2270;
    wire N__2269;
    wire N__2268;
    wire N__2267;
    wire N__2266;
    wire N__2265;
    wire N__2264;
    wire N__2261;
    wire N__2256;
    wire N__2245;
    wire N__2238;
    wire N__2235;
    wire N__2232;
    wire N__2229;
    wire N__2226;
    wire N__2223;
    wire N__2220;
    wire N__2217;
    wire N__2214;
    wire N__2211;
    wire N__2208;
    wire N__2205;
    wire N__2202;
    wire N__2199;
    wire N__2196;
    wire N__2193;
    wire N__2190;
    wire N__2187;
    wire N__2184;
    wire N__2181;
    wire N__2178;
    wire N__2177;
    wire N__2174;
    wire N__2171;
    wire N__2166;
    wire N__2163;
    wire N__2160;
    wire N__2157;
    wire N__2154;
    wire N__2151;
    wire N__2148;
    wire N__2145;
    wire N__2142;
    wire N__2139;
    wire N__2136;
    wire N__2133;
    wire N__2130;
    wire N__2127;
    wire N__2124;
    wire N__2121;
    wire N__2118;
    wire N__2115;
    wire N__2112;
    wire N__2109;
    wire N__2106;
    wire N__2103;
    wire N__2100;
    wire N__2097;
    wire N__2094;
    wire N__2091;
    wire N__2088;
    wire N__2085;
    wire N__2082;
    wire N__2079;
    wire N__2076;
    wire N__2075;
    wire N__2072;
    wire N__2067;
    wire N__2064;
    wire N__2063;
    wire N__2060;
    wire N__2057;
    wire N__2054;
    wire N__2049;
    wire N__2048;
    wire N__2043;
    wire N__2040;
    wire N__2037;
    wire N__2034;
    wire N__2031;
    wire N__2028;
    wire N__2025;
    wire N__2022;
    wire N__2019;
    wire N__2018;
    wire N__2013;
    wire N__2010;
    wire N__2007;
    wire N__2004;
    wire N__2001;
    wire N__1998;
    wire N__1995;
    wire N__1992;
    wire N__1989;
    wire N__1986;
    wire io_jtag_tck_pad_gb_input;
    wire VCCG0;
    wire GNDG0;
    wire n12_cascade_;
    wire n1307;
    wire n2116_cascade_;
    wire n9_adj_2_cascade_;
    wire n8;
    wire n12;
    wire n2_cascade_;
    wire ctrl_idcodeArea_shifter_2;
    wire n1828;
    wire n2045_cascade_;
    wire ctrl_idcodeArea_shifter_4;
    wire ctrl_idcodeArea_shifter_3;
    wire ctrl_idcodeArea_shifter_30;
    wire n1854_cascade_;
    wire n2188_cascade_;
    wire n2235_cascade_;
    wire n2202_cascade_;
    wire n2211;
    wire n962;
    wire n1025;
    wire n1025_cascade_;
    wire n960_cascade_;
    wire n2194;
    wire n1023;
    wire n1027;
    wire n965;
    wire n5;
    wire n5_cascade_;
    wire n2201;
    wire bfn_1_6_0_;
    wire n2009;
    wire n2010;
    wire n2011;
    wire n2012;
    wire n2013;
    wire n2014;
    wire n2015;
    wire n2016;
    wire bfn_1_7_0_;
    wire n2017;
    wire n2018;
    wire n2019;
    wire n2020;
    wire n2021;
    wire n2022;
    wire n2023;
    wire n2024;
    wire bfn_1_8_0_;
    wire n2025;
    wire n2026;
    wire n2027;
    wire n2028;
    wire n2029;
    wire n2030;
    wire n2116;
    wire n4_cascade_;
    wire ctrl_tap_tdoUnbufferd_N_223_cascade_;
    wire ctrl_tap_tdoUnbufferd;
    wire n2146;
    wire n1313_cascade_;
    wire ctrl_tap_tdoUnbufferd_N_224;
    wire ctrl_idcodeArea_shifter_1;
    wire ctrl_idcodeArea_shifter_0;
    wire ctrl_idcodeArea_shifter_29;
    wire ctrl_idcodeArea_shifter_28;
    wire ctrl_idcodeArea_shifter_27;
    wire ctrl_idcodeArea_shifter_26;
    wire ctrl_idcodeArea_shifter_25;
    wire n6;
    wire n1293;
    wire n1582_cascade_;
    wire n2119;
    wire ctrl_idcodeArea_shifter_24;
    wire n2178_cascade_;
    wire ctrl_idcodeArea_shifter_23;
    wire ctrl_idcodeArea_shifter_5;
    wire ctrl_idcodeArea_shifter_7;
    wire ctrl_idcodeArea_shifter_6;
    wire n2045;
    wire ctrl_idcodeArea_shifter_8;
    wire n2140;
    wire n9_cascade_;
    wire n2191;
    wire n12_adj_3;
    wire n1769;
    wire n1864;
    wire myClockArea_timeout_counter_value_3;
    wire myClockArea_timeout_counter_value_1;
    wire myClockArea_timeout_counter_value_5;
    wire myClockArea_timeout_counter_value_0;
    wire myClockArea_timeout_counter_value_9;
    wire myClockArea_timeout_counter_value_18;
    wire myClockArea_timeout_counter_value_12;
    wire myClockArea_timeout_counter_value_14;
    wire ctrl_idcodeArea_shifter_9;
    wire myClockArea_timeout_counter_value_7;
    wire myClockArea_timeout_counter_value_21;
    wire ctrl_idcodeArea_shifter_11;
    wire ctrl_idcodeArea_shifter_10;
    wire myClockArea_timeout_counter_value_4;
    wire myClockArea_timeout_counter_value_6;
    wire myClockArea_timeout_counter_value_22;
    wire myClockArea_timeout_counter_value_16;
    wire myClockArea_timeout_counter_value_17;
    wire myClockArea_timeout_counter_value_8;
    wire myClockArea_timeout_counter_value_10;
    wire myClockArea_timeout_counter_value_2;
    wire n2176;
    wire n2160_cascade_;
    wire n2164;
    wire myClockArea_timeout_counter_value_13;
    wire n11;
    wire n2182_cascade_;
    wire n13;
    wire n2113_cascade_;
    wire n1771;
    wire myClockArea_timeout_counter_value_19;
    wire myClockArea_timeout_counter_value_15;
    wire myClockArea_timeout_counter_value_20;
    wire myClockArea_timeout_counter_value_11;
    wire n2162;
    wire n2113;
    wire global_reset_c;
    wire ctrl_tap_instruction_1;
    wire ctrl_tap_instruction_2;
    wire ctrl_tap_instructionShift_2;
    wire ctrl_tap_instruction_4;
    wire ctrl_tap_instruction_5;
    wire ctrl_tap_instructionShift_5;
    wire ctrl_tap_instruction_7;
    wire ctrl_tap_instructionShift_4;
    wire ctrl_tap_instruction_3;
    wire ctrl_tap_instructionShift_3;
    wire ctrl_tap_instructionShift_7;
    wire ctrl_tap_instruction_6;
    wire ctrl_tap_instructionShift_6;
    wire ctrl_tap_instructionShift_1;
    wire ctrl_tap_instruction_0;
    wire ctrl_tap_instructionShift_0;
    wire n15;
    wire ctrl_idcodeArea_shifter_18;
    wire ctrl_idcodeArea_shifter_20;
    wire ctrl_idcodeArea_shifter_19;
    wire ctrl_idcodeArea_shifter_31;
    wire ctrl_tap_fsm_state_2;
    wire n1067;
    wire ctrl_idcodeArea_shifter_22;
    wire ctrl_idcodeArea_shifter_21;
    wire io_leds_c_0;
    wire ctrl_ledsArea_shifter_0;
    wire io_leds_c_1;
    wire ctrl_ledsArea_shifter_1;
    wire io_leds_c_2;
    wire ctrl_ledsArea_shifter_2;
    wire io_leds_c_3;
    wire ctrl_ledsArea_shifter_3;
    wire ctrl_ledsArea_store_4;
    wire ctrl_ledsArea_shifter_4;
    wire io_leds_c_5;
    wire ctrl_ledsArea_shifter_5;
    wire io_leds_c_6;
    wire ctrl_ledsArea_shifter_6;
    wire n7_adj_1;
    wire io_leds_c_7;
    wire n7;
    wire ctrl_ledsArea_shifter_7;
    wire n1353;
    wire ctrl_tap_fsm_state_0;
    wire ctrl_tap_fsm_state_3;
    wire ctrl_tap_fsm_stateNext_3__N_10_c_3;
    wire ctrl_tap_fsm_state_1;
    wire n963;
    wire myClockArea_timeout_state;
    wire io_leds_c_4;
    wire global_clk_c;
    wire io_jtag_tdi_c;
    wire ctrl_tap_bypass;
    wire ctrl_idcodeArea_shifter_17;
    wire ctrl_idcodeArea_shifter_14;
    wire ctrl_idcodeArea_shifter_13;
    wire ctrl_idcodeArea_shifter_12;
    wire ctrl_idcodeArea_shifter_16;
    wire n2178;
    wire n1582;
    wire ctrl_idcodeArea_shifter_15;
    wire io_jtag_tck_c;
    wire _gnd_net_;

    PRE_IO_GBUF global_clk_pad_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__5398),
            .GLOBALBUFFEROUTPUT(global_clk_c));
    defparam global_clk_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam global_clk_pad_iopad.PULLUP=1'b0;
    IO_PAD global_clk_pad_iopad (
            .OE(N__5400),
            .DIN(N__5399),
            .DOUT(N__5398),
            .PACKAGEPIN(global_clk));
    defparam global_clk_pad_preio.PIN_TYPE=6'b000001;
    defparam global_clk_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO global_clk_pad_preio (
            .PADOEN(N__5400),
            .PADOUT(N__5399),
            .PADIN(N__5398),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam ctrl_tap_fsm_stateNext_3__N_10_pad_3_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ctrl_tap_fsm_stateNext_3__N_10_pad_3_iopad.PULLUP=1'b0;
    IO_PAD ctrl_tap_fsm_stateNext_3__N_10_pad_3_iopad (
            .OE(N__5389),
            .DIN(N__5388),
            .DOUT(N__5387),
            .PACKAGEPIN(io_jtag_tms));
    defparam ctrl_tap_fsm_stateNext_3__N_10_pad_3_preio.PIN_TYPE=6'b000001;
    defparam ctrl_tap_fsm_stateNext_3__N_10_pad_3_preio.NEG_TRIGGER=1'b0;
    PRE_IO ctrl_tap_fsm_stateNext_3__N_10_pad_3_preio (
            .PADOEN(N__5389),
            .PADOUT(N__5388),
            .PADIN(N__5387),
            .CLOCKENABLE(),
            .DIN0(ctrl_tap_fsm_stateNext_3__N_10_c_3),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam global_reset_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam global_reset_pad_iopad.PULLUP=1'b0;
    IO_PAD global_reset_pad_iopad (
            .OE(N__5380),
            .DIN(N__5379),
            .DOUT(N__5378),
            .PACKAGEPIN(global_reset));
    defparam global_reset_pad_preio.PIN_TYPE=6'b000001;
    defparam global_reset_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO global_reset_pad_preio (
            .PADOEN(N__5380),
            .PADOUT(N__5379),
            .PADIN(N__5378),
            .CLOCKENABLE(),
            .DIN0(global_reset_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam io_jtag_tdi_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam io_jtag_tdi_pad_iopad.PULLUP=1'b0;
    IO_PAD io_jtag_tdi_pad_iopad (
            .OE(N__5371),
            .DIN(N__5370),
            .DOUT(N__5369),
            .PACKAGEPIN(io_jtag_tdi));
    defparam io_jtag_tdi_pad_preio.PIN_TYPE=6'b000001;
    defparam io_jtag_tdi_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO io_jtag_tdi_pad_preio (
            .PADOEN(N__5371),
            .PADOUT(N__5370),
            .PADIN(N__5369),
            .CLOCKENABLE(),
            .DIN0(io_jtag_tdi_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam io_jtag_tdo_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam io_jtag_tdo_pad_iopad.PULLUP=1'b0;
    IO_PAD io_jtag_tdo_pad_iopad (
            .OE(N__5362),
            .DIN(N__5361),
            .DOUT(N__5360),
            .PACKAGEPIN(io_jtag_tdo));
    defparam io_jtag_tdo_pad_preio.PIN_TYPE=6'b010101;
    defparam io_jtag_tdo_pad_preio.NEG_TRIGGER=1'b1;
    PRE_IO io_jtag_tdo_pad_preio (
            .PADOEN(N__5362),
            .PADOUT(N__5361),
            .PADIN(N__5360),
            .CLOCKENABLE(VCCG0),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__2283),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(N__4716),
            .OUTPUTENABLE());
    defparam io_leds_pad_0_iopad.IO_STANDARD="SB_LVCMOS";
    defparam io_leds_pad_0_iopad.PULLUP=1'b0;
    IO_PAD io_leds_pad_0_iopad (
            .OE(N__5353),
            .DIN(N__5352),
            .DOUT(N__5351),
            .PACKAGEPIN(io_leds[0]));
    defparam io_leds_pad_0_preio.PIN_TYPE=6'b011001;
    defparam io_leds_pad_0_preio.NEG_TRIGGER=1'b0;
    PRE_IO io_leds_pad_0_preio (
            .PADOEN(N__5353),
            .PADOUT(N__5352),
            .PADIN(N__5351),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__3546),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam io_leds_pad_1_iopad.IO_STANDARD="SB_LVCMOS";
    defparam io_leds_pad_1_iopad.PULLUP=1'b0;
    IO_PAD io_leds_pad_1_iopad (
            .OE(N__5344),
            .DIN(N__5343),
            .DOUT(N__5342),
            .PACKAGEPIN(io_leds[1]));
    defparam io_leds_pad_1_preio.PIN_TYPE=6'b011001;
    defparam io_leds_pad_1_preio.NEG_TRIGGER=1'b0;
    PRE_IO io_leds_pad_1_preio (
            .PADOEN(N__5344),
            .PADOUT(N__5343),
            .PADIN(N__5342),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__4659),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam io_leds_pad_2_iopad.IO_STANDARD="SB_LVCMOS";
    defparam io_leds_pad_2_iopad.PULLUP=1'b0;
    IO_PAD io_leds_pad_2_iopad (
            .OE(N__5335),
            .DIN(N__5334),
            .DOUT(N__5333),
            .PACKAGEPIN(io_leds[2]));
    defparam io_leds_pad_2_preio.PIN_TYPE=6'b011001;
    defparam io_leds_pad_2_preio.NEG_TRIGGER=1'b0;
    PRE_IO io_leds_pad_2_preio (
            .PADOEN(N__5335),
            .PADOUT(N__5334),
            .PADIN(N__5333),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__4605),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam io_leds_pad_3_iopad.IO_STANDARD="SB_LVCMOS";
    defparam io_leds_pad_3_iopad.PULLUP=1'b0;
    IO_PAD io_leds_pad_3_iopad (
            .OE(N__5326),
            .DIN(N__5325),
            .DOUT(N__5324),
            .PACKAGEPIN(io_leds[3]));
    defparam io_leds_pad_3_preio.PIN_TYPE=6'b011001;
    defparam io_leds_pad_3_preio.NEG_TRIGGER=1'b0;
    PRE_IO io_leds_pad_3_preio (
            .PADOEN(N__5326),
            .PADOUT(N__5325),
            .PADIN(N__5324),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__4557),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam io_leds_pad_4_iopad.IO_STANDARD="SB_LVCMOS";
    defparam io_leds_pad_4_iopad.PULLUP=1'b0;
    IO_PAD io_leds_pad_4_iopad (
            .OE(N__5317),
            .DIN(N__5316),
            .DOUT(N__5315),
            .PACKAGEPIN(io_leds[4]));
    defparam io_leds_pad_4_preio.PIN_TYPE=6'b011001;
    defparam io_leds_pad_4_preio.NEG_TRIGGER=1'b0;
    PRE_IO io_leds_pad_4_preio (
            .PADOEN(N__5317),
            .PADOUT(N__5316),
            .PADIN(N__5315),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__5238),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam io_leds_pad_5_iopad.IO_STANDARD="SB_LVCMOS";
    defparam io_leds_pad_5_iopad.PULLUP=1'b0;
    IO_PAD io_leds_pad_5_iopad (
            .OE(N__5308),
            .DIN(N__5307),
            .DOUT(N__5306),
            .PACKAGEPIN(io_leds[5]));
    defparam io_leds_pad_5_preio.PIN_TYPE=6'b011001;
    defparam io_leds_pad_5_preio.NEG_TRIGGER=1'b0;
    PRE_IO io_leds_pad_5_preio (
            .PADOEN(N__5308),
            .PADOUT(N__5307),
            .PADIN(N__5306),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__4464),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam io_leds_pad_6_iopad.IO_STANDARD="SB_LVCMOS";
    defparam io_leds_pad_6_iopad.PULLUP=1'b0;
    IO_PAD io_leds_pad_6_iopad (
            .OE(N__5299),
            .DIN(N__5298),
            .DOUT(N__5297),
            .PACKAGEPIN(io_leds[6]));
    defparam io_leds_pad_6_preio.PIN_TYPE=6'b011001;
    defparam io_leds_pad_6_preio.NEG_TRIGGER=1'b0;
    PRE_IO io_leds_pad_6_preio (
            .PADOEN(N__5299),
            .PADOUT(N__5298),
            .PADIN(N__5297),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__4412),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam io_leds_pad_7_iopad.IO_STANDARD="SB_LVCMOS";
    defparam io_leds_pad_7_iopad.PULLUP=1'b0;
    IO_PAD io_leds_pad_7_iopad (
            .OE(N__5290),
            .DIN(N__5289),
            .DOUT(N__5288),
            .PACKAGEPIN(io_leds[7]));
    defparam io_leds_pad_7_preio.PIN_TYPE=6'b011001;
    defparam io_leds_pad_7_preio.NEG_TRIGGER=1'b0;
    PRE_IO io_leds_pad_7_preio (
            .PADOEN(N__5290),
            .PADOUT(N__5289),
            .PADIN(N__5288),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__4320),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam io_jtag_tck_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam io_jtag_tck_pad_iopad.PULLUP=1'b0;
    IO_PAD io_jtag_tck_pad_iopad (
            .OE(N__5281),
            .DIN(N__5280),
            .DOUT(N__5279),
            .PACKAGEPIN(io_jtag_tck));
    defparam io_jtag_tck_pad_preio.PIN_TYPE=6'b000001;
    defparam io_jtag_tck_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO io_jtag_tck_pad_preio (
            .PADOEN(N__5281),
            .PADOUT(N__5280),
            .PADIN(N__5279),
            .CLOCKENABLE(),
            .DIN0(io_jtag_tck_pad_gb_input),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    InMux I__1261 (
            .O(N__5262),
            .I(N__5258));
    InMux I__1260 (
            .O(N__5261),
            .I(N__5254));
    LocalMux I__1259 (
            .O(N__5258),
            .I(N__5251));
    InMux I__1258 (
            .O(N__5257),
            .I(N__5248));
    LocalMux I__1257 (
            .O(N__5254),
            .I(N__5245));
    Odrv4 I__1256 (
            .O(N__5251),
            .I(myClockArea_timeout_state));
    LocalMux I__1255 (
            .O(N__5248),
            .I(myClockArea_timeout_state));
    Odrv4 I__1254 (
            .O(N__5245),
            .I(myClockArea_timeout_state));
    IoInMux I__1253 (
            .O(N__5238),
            .I(N__5235));
    LocalMux I__1252 (
            .O(N__5235),
            .I(N__5232));
    IoSpan4Mux I__1251 (
            .O(N__5232),
            .I(N__5229));
    Sp12to4 I__1250 (
            .O(N__5229),
            .I(N__5225));
    InMux I__1249 (
            .O(N__5228),
            .I(N__5222));
    Odrv12 I__1248 (
            .O(N__5225),
            .I(io_leds_c_4));
    LocalMux I__1247 (
            .O(N__5222),
            .I(io_leds_c_4));
    ClkMux I__1246 (
            .O(N__5217),
            .I(N__5202));
    ClkMux I__1245 (
            .O(N__5216),
            .I(N__5202));
    ClkMux I__1244 (
            .O(N__5215),
            .I(N__5202));
    ClkMux I__1243 (
            .O(N__5214),
            .I(N__5202));
    ClkMux I__1242 (
            .O(N__5213),
            .I(N__5202));
    GlobalMux I__1241 (
            .O(N__5202),
            .I(N__5199));
    gio2CtrlBuf I__1240 (
            .O(N__5199),
            .I(global_clk_c));
    CascadeMux I__1239 (
            .O(N__5196),
            .I(N__5192));
    CascadeMux I__1238 (
            .O(N__5195),
            .I(N__5189));
    InMux I__1237 (
            .O(N__5192),
            .I(N__5186));
    InMux I__1236 (
            .O(N__5189),
            .I(N__5182));
    LocalMux I__1235 (
            .O(N__5186),
            .I(N__5178));
    InMux I__1234 (
            .O(N__5185),
            .I(N__5175));
    LocalMux I__1233 (
            .O(N__5182),
            .I(N__5172));
    InMux I__1232 (
            .O(N__5181),
            .I(N__5169));
    Span4Mux_v I__1231 (
            .O(N__5178),
            .I(N__5164));
    LocalMux I__1230 (
            .O(N__5175),
            .I(N__5164));
    Odrv4 I__1229 (
            .O(N__5172),
            .I(io_jtag_tdi_c));
    LocalMux I__1228 (
            .O(N__5169),
            .I(io_jtag_tdi_c));
    Odrv4 I__1227 (
            .O(N__5164),
            .I(io_jtag_tdi_c));
    InMux I__1226 (
            .O(N__5157),
            .I(N__5154));
    LocalMux I__1225 (
            .O(N__5154),
            .I(N__5151));
    Odrv4 I__1224 (
            .O(N__5151),
            .I(ctrl_tap_bypass));
    CascadeMux I__1223 (
            .O(N__5148),
            .I(N__5145));
    InMux I__1222 (
            .O(N__5145),
            .I(N__5141));
    InMux I__1221 (
            .O(N__5144),
            .I(N__5138));
    LocalMux I__1220 (
            .O(N__5141),
            .I(ctrl_idcodeArea_shifter_17));
    LocalMux I__1219 (
            .O(N__5138),
            .I(ctrl_idcodeArea_shifter_17));
    InMux I__1218 (
            .O(N__5133),
            .I(N__5127));
    InMux I__1217 (
            .O(N__5132),
            .I(N__5127));
    LocalMux I__1216 (
            .O(N__5127),
            .I(ctrl_idcodeArea_shifter_14));
    CascadeMux I__1215 (
            .O(N__5124),
            .I(N__5121));
    InMux I__1214 (
            .O(N__5121),
            .I(N__5115));
    InMux I__1213 (
            .O(N__5120),
            .I(N__5115));
    LocalMux I__1212 (
            .O(N__5115),
            .I(ctrl_idcodeArea_shifter_13));
    CascadeMux I__1211 (
            .O(N__5112),
            .I(N__5109));
    InMux I__1210 (
            .O(N__5109),
            .I(N__5106));
    LocalMux I__1209 (
            .O(N__5106),
            .I(N__5103));
    Span4Mux_h I__1208 (
            .O(N__5103),
            .I(N__5099));
    InMux I__1207 (
            .O(N__5102),
            .I(N__5096));
    Odrv4 I__1206 (
            .O(N__5099),
            .I(ctrl_idcodeArea_shifter_12));
    LocalMux I__1205 (
            .O(N__5096),
            .I(ctrl_idcodeArea_shifter_12));
    InMux I__1204 (
            .O(N__5091),
            .I(N__5085));
    InMux I__1203 (
            .O(N__5090),
            .I(N__5085));
    LocalMux I__1202 (
            .O(N__5085),
            .I(ctrl_idcodeArea_shifter_16));
    CascadeMux I__1201 (
            .O(N__5082),
            .I(N__5079));
    InMux I__1200 (
            .O(N__5079),
            .I(N__5071));
    InMux I__1199 (
            .O(N__5078),
            .I(N__5068));
    CascadeMux I__1198 (
            .O(N__5077),
            .I(N__5065));
    CascadeMux I__1197 (
            .O(N__5076),
            .I(N__5058));
    InMux I__1196 (
            .O(N__5075),
            .I(N__5032));
    InMux I__1195 (
            .O(N__5074),
            .I(N__5032));
    LocalMux I__1194 (
            .O(N__5071),
            .I(N__5027));
    LocalMux I__1193 (
            .O(N__5068),
            .I(N__5027));
    InMux I__1192 (
            .O(N__5065),
            .I(N__5024));
    InMux I__1191 (
            .O(N__5064),
            .I(N__5021));
    InMux I__1190 (
            .O(N__5063),
            .I(N__5014));
    InMux I__1189 (
            .O(N__5062),
            .I(N__5014));
    InMux I__1188 (
            .O(N__5061),
            .I(N__5014));
    InMux I__1187 (
            .O(N__5058),
            .I(N__5011));
    InMux I__1186 (
            .O(N__5057),
            .I(N__5002));
    InMux I__1185 (
            .O(N__5056),
            .I(N__5002));
    InMux I__1184 (
            .O(N__5055),
            .I(N__5002));
    InMux I__1183 (
            .O(N__5054),
            .I(N__5002));
    InMux I__1182 (
            .O(N__5053),
            .I(N__4991));
    InMux I__1181 (
            .O(N__5052),
            .I(N__4991));
    InMux I__1180 (
            .O(N__5051),
            .I(N__4991));
    InMux I__1179 (
            .O(N__5050),
            .I(N__4991));
    InMux I__1178 (
            .O(N__5049),
            .I(N__4991));
    InMux I__1177 (
            .O(N__5048),
            .I(N__4986));
    InMux I__1176 (
            .O(N__5047),
            .I(N__4986));
    InMux I__1175 (
            .O(N__5046),
            .I(N__4979));
    InMux I__1174 (
            .O(N__5045),
            .I(N__4979));
    InMux I__1173 (
            .O(N__5044),
            .I(N__4979));
    InMux I__1172 (
            .O(N__5043),
            .I(N__4968));
    InMux I__1171 (
            .O(N__5042),
            .I(N__4968));
    InMux I__1170 (
            .O(N__5041),
            .I(N__4968));
    InMux I__1169 (
            .O(N__5040),
            .I(N__4968));
    InMux I__1168 (
            .O(N__5039),
            .I(N__4968));
    InMux I__1167 (
            .O(N__5038),
            .I(N__4963));
    InMux I__1166 (
            .O(N__5037),
            .I(N__4963));
    LocalMux I__1165 (
            .O(N__5032),
            .I(N__4956));
    Span12Mux_s2_v I__1164 (
            .O(N__5027),
            .I(N__4956));
    LocalMux I__1163 (
            .O(N__5024),
            .I(N__4956));
    LocalMux I__1162 (
            .O(N__5021),
            .I(N__4951));
    LocalMux I__1161 (
            .O(N__5014),
            .I(N__4951));
    LocalMux I__1160 (
            .O(N__5011),
            .I(N__4944));
    LocalMux I__1159 (
            .O(N__5002),
            .I(N__4944));
    LocalMux I__1158 (
            .O(N__4991),
            .I(N__4944));
    LocalMux I__1157 (
            .O(N__4986),
            .I(n2178));
    LocalMux I__1156 (
            .O(N__4979),
            .I(n2178));
    LocalMux I__1155 (
            .O(N__4968),
            .I(n2178));
    LocalMux I__1154 (
            .O(N__4963),
            .I(n2178));
    Odrv12 I__1153 (
            .O(N__4956),
            .I(n2178));
    Odrv4 I__1152 (
            .O(N__4951),
            .I(n2178));
    Odrv4 I__1151 (
            .O(N__4944),
            .I(n2178));
    CascadeMux I__1150 (
            .O(N__4929),
            .I(N__4907));
    CascadeMux I__1149 (
            .O(N__4928),
            .I(N__4901));
    InMux I__1148 (
            .O(N__4927),
            .I(N__4885));
    InMux I__1147 (
            .O(N__4926),
            .I(N__4885));
    InMux I__1146 (
            .O(N__4925),
            .I(N__4885));
    InMux I__1145 (
            .O(N__4924),
            .I(N__4885));
    InMux I__1144 (
            .O(N__4923),
            .I(N__4885));
    InMux I__1143 (
            .O(N__4922),
            .I(N__4878));
    InMux I__1142 (
            .O(N__4921),
            .I(N__4878));
    InMux I__1141 (
            .O(N__4920),
            .I(N__4878));
    CascadeMux I__1140 (
            .O(N__4919),
            .I(N__4874));
    CascadeMux I__1139 (
            .O(N__4918),
            .I(N__4871));
    CascadeMux I__1138 (
            .O(N__4917),
            .I(N__4867));
    CascadeMux I__1137 (
            .O(N__4916),
            .I(N__4860));
    InMux I__1136 (
            .O(N__4915),
            .I(N__4851));
    InMux I__1135 (
            .O(N__4914),
            .I(N__4848));
    InMux I__1134 (
            .O(N__4913),
            .I(N__4841));
    InMux I__1133 (
            .O(N__4912),
            .I(N__4841));
    InMux I__1132 (
            .O(N__4911),
            .I(N__4841));
    InMux I__1131 (
            .O(N__4910),
            .I(N__4832));
    InMux I__1130 (
            .O(N__4907),
            .I(N__4832));
    InMux I__1129 (
            .O(N__4906),
            .I(N__4832));
    InMux I__1128 (
            .O(N__4905),
            .I(N__4832));
    InMux I__1127 (
            .O(N__4904),
            .I(N__4825));
    InMux I__1126 (
            .O(N__4901),
            .I(N__4825));
    InMux I__1125 (
            .O(N__4900),
            .I(N__4825));
    InMux I__1124 (
            .O(N__4899),
            .I(N__4822));
    InMux I__1123 (
            .O(N__4898),
            .I(N__4815));
    InMux I__1122 (
            .O(N__4897),
            .I(N__4815));
    InMux I__1121 (
            .O(N__4896),
            .I(N__4815));
    LocalMux I__1120 (
            .O(N__4885),
            .I(N__4810));
    LocalMux I__1119 (
            .O(N__4878),
            .I(N__4810));
    InMux I__1118 (
            .O(N__4877),
            .I(N__4807));
    InMux I__1117 (
            .O(N__4874),
            .I(N__4804));
    InMux I__1116 (
            .O(N__4871),
            .I(N__4801));
    InMux I__1115 (
            .O(N__4870),
            .I(N__4796));
    InMux I__1114 (
            .O(N__4867),
            .I(N__4796));
    InMux I__1113 (
            .O(N__4866),
            .I(N__4791));
    InMux I__1112 (
            .O(N__4865),
            .I(N__4791));
    InMux I__1111 (
            .O(N__4864),
            .I(N__4786));
    InMux I__1110 (
            .O(N__4863),
            .I(N__4786));
    InMux I__1109 (
            .O(N__4860),
            .I(N__4779));
    InMux I__1108 (
            .O(N__4859),
            .I(N__4779));
    InMux I__1107 (
            .O(N__4858),
            .I(N__4779));
    InMux I__1106 (
            .O(N__4857),
            .I(N__4770));
    InMux I__1105 (
            .O(N__4856),
            .I(N__4770));
    InMux I__1104 (
            .O(N__4855),
            .I(N__4770));
    InMux I__1103 (
            .O(N__4854),
            .I(N__4770));
    LocalMux I__1102 (
            .O(N__4851),
            .I(N__4767));
    LocalMux I__1101 (
            .O(N__4848),
            .I(N__4758));
    LocalMux I__1100 (
            .O(N__4841),
            .I(N__4758));
    LocalMux I__1099 (
            .O(N__4832),
            .I(N__4758));
    LocalMux I__1098 (
            .O(N__4825),
            .I(N__4758));
    LocalMux I__1097 (
            .O(N__4822),
            .I(N__4751));
    LocalMux I__1096 (
            .O(N__4815),
            .I(N__4751));
    Span4Mux_s1_v I__1095 (
            .O(N__4810),
            .I(N__4751));
    LocalMux I__1094 (
            .O(N__4807),
            .I(n1582));
    LocalMux I__1093 (
            .O(N__4804),
            .I(n1582));
    LocalMux I__1092 (
            .O(N__4801),
            .I(n1582));
    LocalMux I__1091 (
            .O(N__4796),
            .I(n1582));
    LocalMux I__1090 (
            .O(N__4791),
            .I(n1582));
    LocalMux I__1089 (
            .O(N__4786),
            .I(n1582));
    LocalMux I__1088 (
            .O(N__4779),
            .I(n1582));
    LocalMux I__1087 (
            .O(N__4770),
            .I(n1582));
    Odrv4 I__1086 (
            .O(N__4767),
            .I(n1582));
    Odrv4 I__1085 (
            .O(N__4758),
            .I(n1582));
    Odrv4 I__1084 (
            .O(N__4751),
            .I(n1582));
    CascadeMux I__1083 (
            .O(N__4728),
            .I(N__4724));
    InMux I__1082 (
            .O(N__4727),
            .I(N__4719));
    InMux I__1081 (
            .O(N__4724),
            .I(N__4719));
    LocalMux I__1080 (
            .O(N__4719),
            .I(ctrl_idcodeArea_shifter_15));
    ClkMux I__1079 (
            .O(N__4716),
            .I(N__4665));
    ClkMux I__1078 (
            .O(N__4715),
            .I(N__4665));
    ClkMux I__1077 (
            .O(N__4714),
            .I(N__4665));
    ClkMux I__1076 (
            .O(N__4713),
            .I(N__4665));
    ClkMux I__1075 (
            .O(N__4712),
            .I(N__4665));
    ClkMux I__1074 (
            .O(N__4711),
            .I(N__4665));
    ClkMux I__1073 (
            .O(N__4710),
            .I(N__4665));
    ClkMux I__1072 (
            .O(N__4709),
            .I(N__4665));
    ClkMux I__1071 (
            .O(N__4708),
            .I(N__4665));
    ClkMux I__1070 (
            .O(N__4707),
            .I(N__4665));
    ClkMux I__1069 (
            .O(N__4706),
            .I(N__4665));
    ClkMux I__1068 (
            .O(N__4705),
            .I(N__4665));
    ClkMux I__1067 (
            .O(N__4704),
            .I(N__4665));
    ClkMux I__1066 (
            .O(N__4703),
            .I(N__4665));
    ClkMux I__1065 (
            .O(N__4702),
            .I(N__4665));
    ClkMux I__1064 (
            .O(N__4701),
            .I(N__4665));
    ClkMux I__1063 (
            .O(N__4700),
            .I(N__4665));
    GlobalMux I__1062 (
            .O(N__4665),
            .I(N__4662));
    gio2CtrlBuf I__1061 (
            .O(N__4662),
            .I(io_jtag_tck_c));
    IoInMux I__1060 (
            .O(N__4659),
            .I(N__4656));
    LocalMux I__1059 (
            .O(N__4656),
            .I(N__4653));
    Span4Mux_s2_h I__1058 (
            .O(N__4653),
            .I(N__4650));
    Span4Mux_h I__1057 (
            .O(N__4650),
            .I(N__4646));
    CascadeMux I__1056 (
            .O(N__4649),
            .I(N__4643));
    Span4Mux_v I__1055 (
            .O(N__4646),
            .I(N__4640));
    InMux I__1054 (
            .O(N__4643),
            .I(N__4637));
    Span4Mux_v I__1053 (
            .O(N__4640),
            .I(N__4631));
    LocalMux I__1052 (
            .O(N__4637),
            .I(N__4631));
    InMux I__1051 (
            .O(N__4636),
            .I(N__4628));
    Odrv4 I__1050 (
            .O(N__4631),
            .I(io_leds_c_1));
    LocalMux I__1049 (
            .O(N__4628),
            .I(io_leds_c_1));
    InMux I__1048 (
            .O(N__4623),
            .I(N__4619));
    CascadeMux I__1047 (
            .O(N__4622),
            .I(N__4616));
    LocalMux I__1046 (
            .O(N__4619),
            .I(N__4613));
    InMux I__1045 (
            .O(N__4616),
            .I(N__4610));
    Odrv4 I__1044 (
            .O(N__4613),
            .I(ctrl_ledsArea_shifter_1));
    LocalMux I__1043 (
            .O(N__4610),
            .I(ctrl_ledsArea_shifter_1));
    IoInMux I__1042 (
            .O(N__4605),
            .I(N__4602));
    LocalMux I__1041 (
            .O(N__4602),
            .I(N__4599));
    Span4Mux_s3_h I__1040 (
            .O(N__4599),
            .I(N__4596));
    Sp12to4 I__1039 (
            .O(N__4596),
            .I(N__4592));
    InMux I__1038 (
            .O(N__4595),
            .I(N__4589));
    Span12Mux_v I__1037 (
            .O(N__4592),
            .I(N__4583));
    LocalMux I__1036 (
            .O(N__4589),
            .I(N__4583));
    InMux I__1035 (
            .O(N__4588),
            .I(N__4580));
    Odrv12 I__1034 (
            .O(N__4583),
            .I(io_leds_c_2));
    LocalMux I__1033 (
            .O(N__4580),
            .I(io_leds_c_2));
    InMux I__1032 (
            .O(N__4575),
            .I(N__4572));
    LocalMux I__1031 (
            .O(N__4572),
            .I(N__4568));
    InMux I__1030 (
            .O(N__4571),
            .I(N__4565));
    Span4Mux_s2_h I__1029 (
            .O(N__4568),
            .I(N__4560));
    LocalMux I__1028 (
            .O(N__4565),
            .I(N__4560));
    Odrv4 I__1027 (
            .O(N__4560),
            .I(ctrl_ledsArea_shifter_2));
    IoInMux I__1026 (
            .O(N__4557),
            .I(N__4554));
    LocalMux I__1025 (
            .O(N__4554),
            .I(N__4551));
    IoSpan4Mux I__1024 (
            .O(N__4551),
            .I(N__4548));
    Span4Mux_s3_h I__1023 (
            .O(N__4548),
            .I(N__4545));
    Span4Mux_h I__1022 (
            .O(N__4545),
            .I(N__4541));
    InMux I__1021 (
            .O(N__4544),
            .I(N__4538));
    Span4Mux_v I__1020 (
            .O(N__4541),
            .I(N__4532));
    LocalMux I__1019 (
            .O(N__4538),
            .I(N__4532));
    InMux I__1018 (
            .O(N__4537),
            .I(N__4529));
    Odrv4 I__1017 (
            .O(N__4532),
            .I(io_leds_c_3));
    LocalMux I__1016 (
            .O(N__4529),
            .I(io_leds_c_3));
    CascadeMux I__1015 (
            .O(N__4524),
            .I(N__4521));
    InMux I__1014 (
            .O(N__4521),
            .I(N__4517));
    CascadeMux I__1013 (
            .O(N__4520),
            .I(N__4514));
    LocalMux I__1012 (
            .O(N__4517),
            .I(N__4511));
    InMux I__1011 (
            .O(N__4514),
            .I(N__4508));
    Odrv4 I__1010 (
            .O(N__4511),
            .I(ctrl_ledsArea_shifter_3));
    LocalMux I__1009 (
            .O(N__4508),
            .I(ctrl_ledsArea_shifter_3));
    InMux I__1008 (
            .O(N__4503),
            .I(N__4500));
    LocalMux I__1007 (
            .O(N__4500),
            .I(N__4497));
    Span4Mux_h I__1006 (
            .O(N__4497),
            .I(N__4493));
    InMux I__1005 (
            .O(N__4496),
            .I(N__4490));
    Odrv4 I__1004 (
            .O(N__4493),
            .I(ctrl_ledsArea_store_4));
    LocalMux I__1003 (
            .O(N__4490),
            .I(ctrl_ledsArea_store_4));
    InMux I__1002 (
            .O(N__4485),
            .I(N__4482));
    LocalMux I__1001 (
            .O(N__4482),
            .I(N__4478));
    CascadeMux I__1000 (
            .O(N__4481),
            .I(N__4475));
    Span4Mux_s3_h I__999 (
            .O(N__4478),
            .I(N__4472));
    InMux I__998 (
            .O(N__4475),
            .I(N__4469));
    Odrv4 I__997 (
            .O(N__4472),
            .I(ctrl_ledsArea_shifter_4));
    LocalMux I__996 (
            .O(N__4469),
            .I(ctrl_ledsArea_shifter_4));
    IoInMux I__995 (
            .O(N__4464),
            .I(N__4461));
    LocalMux I__994 (
            .O(N__4461),
            .I(N__4458));
    Span4Mux_s1_h I__993 (
            .O(N__4458),
            .I(N__4454));
    InMux I__992 (
            .O(N__4457),
            .I(N__4451));
    Span4Mux_v I__991 (
            .O(N__4454),
            .I(N__4447));
    LocalMux I__990 (
            .O(N__4451),
            .I(N__4444));
    InMux I__989 (
            .O(N__4450),
            .I(N__4441));
    Odrv4 I__988 (
            .O(N__4447),
            .I(io_leds_c_5));
    Odrv12 I__987 (
            .O(N__4444),
            .I(io_leds_c_5));
    LocalMux I__986 (
            .O(N__4441),
            .I(io_leds_c_5));
    CascadeMux I__985 (
            .O(N__4434),
            .I(N__4431));
    InMux I__984 (
            .O(N__4431),
            .I(N__4428));
    LocalMux I__983 (
            .O(N__4428),
            .I(N__4424));
    InMux I__982 (
            .O(N__4427),
            .I(N__4421));
    Odrv4 I__981 (
            .O(N__4424),
            .I(ctrl_ledsArea_shifter_5));
    LocalMux I__980 (
            .O(N__4421),
            .I(ctrl_ledsArea_shifter_5));
    InMux I__979 (
            .O(N__4416),
            .I(N__4413));
    LocalMux I__978 (
            .O(N__4413),
            .I(N__4409));
    IoInMux I__977 (
            .O(N__4412),
            .I(N__4405));
    Span4Mux_h I__976 (
            .O(N__4409),
            .I(N__4402));
    InMux I__975 (
            .O(N__4408),
            .I(N__4399));
    LocalMux I__974 (
            .O(N__4405),
            .I(io_leds_c_6));
    Odrv4 I__973 (
            .O(N__4402),
            .I(io_leds_c_6));
    LocalMux I__972 (
            .O(N__4399),
            .I(io_leds_c_6));
    InMux I__971 (
            .O(N__4392),
            .I(N__4389));
    LocalMux I__970 (
            .O(N__4389),
            .I(N__4385));
    CascadeMux I__969 (
            .O(N__4388),
            .I(N__4382));
    Span4Mux_s3_h I__968 (
            .O(N__4385),
            .I(N__4379));
    InMux I__967 (
            .O(N__4382),
            .I(N__4376));
    Odrv4 I__966 (
            .O(N__4379),
            .I(ctrl_ledsArea_shifter_6));
    LocalMux I__965 (
            .O(N__4376),
            .I(ctrl_ledsArea_shifter_6));
    CascadeMux I__964 (
            .O(N__4371),
            .I(N__4368));
    InMux I__963 (
            .O(N__4368),
            .I(N__4358));
    InMux I__962 (
            .O(N__4367),
            .I(N__4343));
    InMux I__961 (
            .O(N__4366),
            .I(N__4343));
    InMux I__960 (
            .O(N__4365),
            .I(N__4343));
    InMux I__959 (
            .O(N__4364),
            .I(N__4343));
    InMux I__958 (
            .O(N__4363),
            .I(N__4343));
    InMux I__957 (
            .O(N__4362),
            .I(N__4343));
    InMux I__956 (
            .O(N__4361),
            .I(N__4343));
    LocalMux I__955 (
            .O(N__4358),
            .I(N__4338));
    LocalMux I__954 (
            .O(N__4343),
            .I(N__4335));
    InMux I__953 (
            .O(N__4342),
            .I(N__4330));
    InMux I__952 (
            .O(N__4341),
            .I(N__4330));
    Span4Mux_h I__951 (
            .O(N__4338),
            .I(N__4323));
    Span4Mux_h I__950 (
            .O(N__4335),
            .I(N__4323));
    LocalMux I__949 (
            .O(N__4330),
            .I(N__4323));
    Odrv4 I__948 (
            .O(N__4323),
            .I(n7_adj_1));
    IoInMux I__947 (
            .O(N__4320),
            .I(N__4317));
    LocalMux I__946 (
            .O(N__4317),
            .I(N__4314));
    Span4Mux_s0_h I__945 (
            .O(N__4314),
            .I(N__4310));
    InMux I__944 (
            .O(N__4313),
            .I(N__4307));
    Span4Mux_v I__943 (
            .O(N__4310),
            .I(N__4303));
    LocalMux I__942 (
            .O(N__4307),
            .I(N__4300));
    InMux I__941 (
            .O(N__4306),
            .I(N__4297));
    Odrv4 I__940 (
            .O(N__4303),
            .I(io_leds_c_7));
    Odrv12 I__939 (
            .O(N__4300),
            .I(io_leds_c_7));
    LocalMux I__938 (
            .O(N__4297),
            .I(io_leds_c_7));
    InMux I__937 (
            .O(N__4290),
            .I(N__4274));
    InMux I__936 (
            .O(N__4289),
            .I(N__4274));
    InMux I__935 (
            .O(N__4288),
            .I(N__4274));
    InMux I__934 (
            .O(N__4287),
            .I(N__4274));
    InMux I__933 (
            .O(N__4286),
            .I(N__4265));
    InMux I__932 (
            .O(N__4285),
            .I(N__4265));
    InMux I__931 (
            .O(N__4284),
            .I(N__4265));
    InMux I__930 (
            .O(N__4283),
            .I(N__4265));
    LocalMux I__929 (
            .O(N__4274),
            .I(N__4260));
    LocalMux I__928 (
            .O(N__4265),
            .I(N__4260));
    Span4Mux_h I__927 (
            .O(N__4260),
            .I(N__4257));
    Odrv4 I__926 (
            .O(N__4257),
            .I(n7));
    InMux I__925 (
            .O(N__4254),
            .I(N__4250));
    CascadeMux I__924 (
            .O(N__4253),
            .I(N__4247));
    LocalMux I__923 (
            .O(N__4250),
            .I(N__4244));
    InMux I__922 (
            .O(N__4247),
            .I(N__4241));
    Odrv4 I__921 (
            .O(N__4244),
            .I(ctrl_ledsArea_shifter_7));
    LocalMux I__920 (
            .O(N__4241),
            .I(ctrl_ledsArea_shifter_7));
    CEMux I__919 (
            .O(N__4236),
            .I(N__4233));
    LocalMux I__918 (
            .O(N__4233),
            .I(N__4230));
    Span4Mux_h I__917 (
            .O(N__4230),
            .I(N__4227));
    Odrv4 I__916 (
            .O(N__4227),
            .I(n1353));
    InMux I__915 (
            .O(N__4224),
            .I(N__4210));
    InMux I__914 (
            .O(N__4223),
            .I(N__4195));
    InMux I__913 (
            .O(N__4222),
            .I(N__4195));
    InMux I__912 (
            .O(N__4221),
            .I(N__4195));
    InMux I__911 (
            .O(N__4220),
            .I(N__4195));
    InMux I__910 (
            .O(N__4219),
            .I(N__4195));
    InMux I__909 (
            .O(N__4218),
            .I(N__4195));
    InMux I__908 (
            .O(N__4217),
            .I(N__4195));
    InMux I__907 (
            .O(N__4216),
            .I(N__4192));
    InMux I__906 (
            .O(N__4215),
            .I(N__4189));
    CascadeMux I__905 (
            .O(N__4214),
            .I(N__4185));
    CascadeMux I__904 (
            .O(N__4213),
            .I(N__4179));
    LocalMux I__903 (
            .O(N__4210),
            .I(N__4161));
    LocalMux I__902 (
            .O(N__4195),
            .I(N__4161));
    LocalMux I__901 (
            .O(N__4192),
            .I(N__4161));
    LocalMux I__900 (
            .O(N__4189),
            .I(N__4158));
    InMux I__899 (
            .O(N__4188),
            .I(N__4151));
    InMux I__898 (
            .O(N__4185),
            .I(N__4151));
    InMux I__897 (
            .O(N__4184),
            .I(N__4151));
    InMux I__896 (
            .O(N__4183),
            .I(N__4148));
    InMux I__895 (
            .O(N__4182),
            .I(N__4141));
    InMux I__894 (
            .O(N__4179),
            .I(N__4141));
    InMux I__893 (
            .O(N__4178),
            .I(N__4138));
    InMux I__892 (
            .O(N__4177),
            .I(N__4127));
    InMux I__891 (
            .O(N__4176),
            .I(N__4127));
    InMux I__890 (
            .O(N__4175),
            .I(N__4127));
    InMux I__889 (
            .O(N__4174),
            .I(N__4127));
    InMux I__888 (
            .O(N__4173),
            .I(N__4127));
    InMux I__887 (
            .O(N__4172),
            .I(N__4116));
    InMux I__886 (
            .O(N__4171),
            .I(N__4116));
    InMux I__885 (
            .O(N__4170),
            .I(N__4116));
    InMux I__884 (
            .O(N__4169),
            .I(N__4116));
    InMux I__883 (
            .O(N__4168),
            .I(N__4116));
    Span4Mux_s3_v I__882 (
            .O(N__4161),
            .I(N__4111));
    Span4Mux_v I__881 (
            .O(N__4158),
            .I(N__4111));
    LocalMux I__880 (
            .O(N__4151),
            .I(N__4106));
    LocalMux I__879 (
            .O(N__4148),
            .I(N__4106));
    InMux I__878 (
            .O(N__4147),
            .I(N__4101));
    InMux I__877 (
            .O(N__4146),
            .I(N__4101));
    LocalMux I__876 (
            .O(N__4141),
            .I(ctrl_tap_fsm_state_0));
    LocalMux I__875 (
            .O(N__4138),
            .I(ctrl_tap_fsm_state_0));
    LocalMux I__874 (
            .O(N__4127),
            .I(ctrl_tap_fsm_state_0));
    LocalMux I__873 (
            .O(N__4116),
            .I(ctrl_tap_fsm_state_0));
    Odrv4 I__872 (
            .O(N__4111),
            .I(ctrl_tap_fsm_state_0));
    Odrv4 I__871 (
            .O(N__4106),
            .I(ctrl_tap_fsm_state_0));
    LocalMux I__870 (
            .O(N__4101),
            .I(ctrl_tap_fsm_state_0));
    InMux I__869 (
            .O(N__4086),
            .I(N__4080));
    InMux I__868 (
            .O(N__4085),
            .I(N__4077));
    InMux I__867 (
            .O(N__4084),
            .I(N__4073));
    CascadeMux I__866 (
            .O(N__4083),
            .I(N__4059));
    LocalMux I__865 (
            .O(N__4080),
            .I(N__4054));
    LocalMux I__864 (
            .O(N__4077),
            .I(N__4054));
    InMux I__863 (
            .O(N__4076),
            .I(N__4048));
    LocalMux I__862 (
            .O(N__4073),
            .I(N__4045));
    InMux I__861 (
            .O(N__4072),
            .I(N__4042));
    CascadeMux I__860 (
            .O(N__4071),
            .I(N__4039));
    InMux I__859 (
            .O(N__4070),
            .I(N__4033));
    InMux I__858 (
            .O(N__4069),
            .I(N__4033));
    InMux I__857 (
            .O(N__4068),
            .I(N__4030));
    InMux I__856 (
            .O(N__4067),
            .I(N__4023));
    InMux I__855 (
            .O(N__4066),
            .I(N__4023));
    InMux I__854 (
            .O(N__4065),
            .I(N__4023));
    InMux I__853 (
            .O(N__4064),
            .I(N__4014));
    InMux I__852 (
            .O(N__4063),
            .I(N__4014));
    InMux I__851 (
            .O(N__4062),
            .I(N__4014));
    InMux I__850 (
            .O(N__4059),
            .I(N__4014));
    Span4Mux_h I__849 (
            .O(N__4054),
            .I(N__4011));
    InMux I__848 (
            .O(N__4053),
            .I(N__4004));
    InMux I__847 (
            .O(N__4052),
            .I(N__4004));
    InMux I__846 (
            .O(N__4051),
            .I(N__4004));
    LocalMux I__845 (
            .O(N__4048),
            .I(N__3997));
    Span4Mux_h I__844 (
            .O(N__4045),
            .I(N__3997));
    LocalMux I__843 (
            .O(N__4042),
            .I(N__3997));
    InMux I__842 (
            .O(N__4039),
            .I(N__3992));
    InMux I__841 (
            .O(N__4038),
            .I(N__3992));
    LocalMux I__840 (
            .O(N__4033),
            .I(ctrl_tap_fsm_state_3));
    LocalMux I__839 (
            .O(N__4030),
            .I(ctrl_tap_fsm_state_3));
    LocalMux I__838 (
            .O(N__4023),
            .I(ctrl_tap_fsm_state_3));
    LocalMux I__837 (
            .O(N__4014),
            .I(ctrl_tap_fsm_state_3));
    Odrv4 I__836 (
            .O(N__4011),
            .I(ctrl_tap_fsm_state_3));
    LocalMux I__835 (
            .O(N__4004),
            .I(ctrl_tap_fsm_state_3));
    Odrv4 I__834 (
            .O(N__3997),
            .I(ctrl_tap_fsm_state_3));
    LocalMux I__833 (
            .O(N__3992),
            .I(ctrl_tap_fsm_state_3));
    CascadeMux I__832 (
            .O(N__3975),
            .I(N__3969));
    CascadeMux I__831 (
            .O(N__3974),
            .I(N__3965));
    CascadeMux I__830 (
            .O(N__3973),
            .I(N__3958));
    InMux I__829 (
            .O(N__3972),
            .I(N__3955));
    InMux I__828 (
            .O(N__3969),
            .I(N__3950));
    InMux I__827 (
            .O(N__3968),
            .I(N__3950));
    InMux I__826 (
            .O(N__3965),
            .I(N__3945));
    InMux I__825 (
            .O(N__3964),
            .I(N__3945));
    InMux I__824 (
            .O(N__3963),
            .I(N__3938));
    InMux I__823 (
            .O(N__3962),
            .I(N__3938));
    InMux I__822 (
            .O(N__3961),
            .I(N__3938));
    InMux I__821 (
            .O(N__3958),
            .I(N__3934));
    LocalMux I__820 (
            .O(N__3955),
            .I(N__3930));
    LocalMux I__819 (
            .O(N__3950),
            .I(N__3923));
    LocalMux I__818 (
            .O(N__3945),
            .I(N__3923));
    LocalMux I__817 (
            .O(N__3938),
            .I(N__3923));
    InMux I__816 (
            .O(N__3937),
            .I(N__3920));
    LocalMux I__815 (
            .O(N__3934),
            .I(N__3917));
    CascadeMux I__814 (
            .O(N__3933),
            .I(N__3914));
    Span4Mux_v I__813 (
            .O(N__3930),
            .I(N__3909));
    Span4Mux_v I__812 (
            .O(N__3923),
            .I(N__3909));
    LocalMux I__811 (
            .O(N__3920),
            .I(N__3906));
    Span4Mux_s3_h I__810 (
            .O(N__3917),
            .I(N__3903));
    InMux I__809 (
            .O(N__3914),
            .I(N__3900));
    IoSpan4Mux I__808 (
            .O(N__3909),
            .I(N__3897));
    Span4Mux_s3_h I__807 (
            .O(N__3906),
            .I(N__3894));
    Sp12to4 I__806 (
            .O(N__3903),
            .I(N__3889));
    LocalMux I__805 (
            .O(N__3900),
            .I(N__3889));
    Odrv4 I__804 (
            .O(N__3897),
            .I(ctrl_tap_fsm_stateNext_3__N_10_c_3));
    Odrv4 I__803 (
            .O(N__3894),
            .I(ctrl_tap_fsm_stateNext_3__N_10_c_3));
    Odrv12 I__802 (
            .O(N__3889),
            .I(ctrl_tap_fsm_stateNext_3__N_10_c_3));
    InMux I__801 (
            .O(N__3882),
            .I(N__3875));
    InMux I__800 (
            .O(N__3881),
            .I(N__3875));
    InMux I__799 (
            .O(N__3880),
            .I(N__3872));
    LocalMux I__798 (
            .O(N__3875),
            .I(N__3865));
    LocalMux I__797 (
            .O(N__3872),
            .I(N__3850));
    InMux I__796 (
            .O(N__3871),
            .I(N__3843));
    InMux I__795 (
            .O(N__3870),
            .I(N__3843));
    InMux I__794 (
            .O(N__3869),
            .I(N__3843));
    InMux I__793 (
            .O(N__3868),
            .I(N__3840));
    Span4Mux_h I__792 (
            .O(N__3865),
            .I(N__3835));
    InMux I__791 (
            .O(N__3864),
            .I(N__3832));
    InMux I__790 (
            .O(N__3863),
            .I(N__3829));
    InMux I__789 (
            .O(N__3862),
            .I(N__3818));
    InMux I__788 (
            .O(N__3861),
            .I(N__3818));
    InMux I__787 (
            .O(N__3860),
            .I(N__3818));
    InMux I__786 (
            .O(N__3859),
            .I(N__3818));
    InMux I__785 (
            .O(N__3858),
            .I(N__3818));
    InMux I__784 (
            .O(N__3857),
            .I(N__3807));
    InMux I__783 (
            .O(N__3856),
            .I(N__3807));
    InMux I__782 (
            .O(N__3855),
            .I(N__3807));
    InMux I__781 (
            .O(N__3854),
            .I(N__3807));
    InMux I__780 (
            .O(N__3853),
            .I(N__3807));
    Span4Mux_h I__779 (
            .O(N__3850),
            .I(N__3800));
    LocalMux I__778 (
            .O(N__3843),
            .I(N__3800));
    LocalMux I__777 (
            .O(N__3840),
            .I(N__3800));
    InMux I__776 (
            .O(N__3839),
            .I(N__3795));
    InMux I__775 (
            .O(N__3838),
            .I(N__3795));
    Odrv4 I__774 (
            .O(N__3835),
            .I(ctrl_tap_fsm_state_1));
    LocalMux I__773 (
            .O(N__3832),
            .I(ctrl_tap_fsm_state_1));
    LocalMux I__772 (
            .O(N__3829),
            .I(ctrl_tap_fsm_state_1));
    LocalMux I__771 (
            .O(N__3818),
            .I(ctrl_tap_fsm_state_1));
    LocalMux I__770 (
            .O(N__3807),
            .I(ctrl_tap_fsm_state_1));
    Odrv4 I__769 (
            .O(N__3800),
            .I(ctrl_tap_fsm_state_1));
    LocalMux I__768 (
            .O(N__3795),
            .I(ctrl_tap_fsm_state_1));
    InMux I__767 (
            .O(N__3780),
            .I(N__3777));
    LocalMux I__766 (
            .O(N__3777),
            .I(N__3774));
    Span4Mux_s3_h I__765 (
            .O(N__3774),
            .I(N__3771));
    Odrv4 I__764 (
            .O(N__3771),
            .I(n963));
    InMux I__763 (
            .O(N__3768),
            .I(N__3765));
    LocalMux I__762 (
            .O(N__3765),
            .I(N__3762));
    Span4Mux_h I__761 (
            .O(N__3762),
            .I(N__3758));
    InMux I__760 (
            .O(N__3761),
            .I(N__3755));
    Odrv4 I__759 (
            .O(N__3758),
            .I(n15));
    LocalMux I__758 (
            .O(N__3755),
            .I(n15));
    CascadeMux I__757 (
            .O(N__3750),
            .I(N__3747));
    InMux I__756 (
            .O(N__3747),
            .I(N__3741));
    InMux I__755 (
            .O(N__3746),
            .I(N__3741));
    LocalMux I__754 (
            .O(N__3741),
            .I(ctrl_idcodeArea_shifter_18));
    CascadeMux I__753 (
            .O(N__3738),
            .I(N__3734));
    InMux I__752 (
            .O(N__3737),
            .I(N__3729));
    InMux I__751 (
            .O(N__3734),
            .I(N__3729));
    LocalMux I__750 (
            .O(N__3729),
            .I(ctrl_idcodeArea_shifter_20));
    InMux I__749 (
            .O(N__3726),
            .I(N__3720));
    InMux I__748 (
            .O(N__3725),
            .I(N__3720));
    LocalMux I__747 (
            .O(N__3720),
            .I(ctrl_idcodeArea_shifter_19));
    InMux I__746 (
            .O(N__3717),
            .I(N__3713));
    InMux I__745 (
            .O(N__3716),
            .I(N__3710));
    LocalMux I__744 (
            .O(N__3713),
            .I(N__3707));
    LocalMux I__743 (
            .O(N__3710),
            .I(ctrl_idcodeArea_shifter_31));
    Odrv12 I__742 (
            .O(N__3707),
            .I(ctrl_idcodeArea_shifter_31));
    CascadeMux I__741 (
            .O(N__3702),
            .I(N__3698));
    CascadeMux I__740 (
            .O(N__3701),
            .I(N__3695));
    InMux I__739 (
            .O(N__3698),
            .I(N__3685));
    InMux I__738 (
            .O(N__3695),
            .I(N__3685));
    CascadeMux I__737 (
            .O(N__3694),
            .I(N__3678));
    CascadeMux I__736 (
            .O(N__3693),
            .I(N__3674));
    CascadeMux I__735 (
            .O(N__3692),
            .I(N__3671));
    CascadeMux I__734 (
            .O(N__3691),
            .I(N__3667));
    CascadeMux I__733 (
            .O(N__3690),
            .I(N__3664));
    LocalMux I__732 (
            .O(N__3685),
            .I(N__3660));
    InMux I__731 (
            .O(N__3684),
            .I(N__3653));
    InMux I__730 (
            .O(N__3683),
            .I(N__3653));
    InMux I__729 (
            .O(N__3682),
            .I(N__3650));
    CascadeMux I__728 (
            .O(N__3681),
            .I(N__3646));
    InMux I__727 (
            .O(N__3678),
            .I(N__3641));
    InMux I__726 (
            .O(N__3677),
            .I(N__3641));
    InMux I__725 (
            .O(N__3674),
            .I(N__3636));
    InMux I__724 (
            .O(N__3671),
            .I(N__3636));
    InMux I__723 (
            .O(N__3670),
            .I(N__3627));
    InMux I__722 (
            .O(N__3667),
            .I(N__3627));
    InMux I__721 (
            .O(N__3664),
            .I(N__3627));
    InMux I__720 (
            .O(N__3663),
            .I(N__3627));
    Span4Mux_h I__719 (
            .O(N__3660),
            .I(N__3624));
    InMux I__718 (
            .O(N__3659),
            .I(N__3619));
    InMux I__717 (
            .O(N__3658),
            .I(N__3619));
    LocalMux I__716 (
            .O(N__3653),
            .I(N__3614));
    LocalMux I__715 (
            .O(N__3650),
            .I(N__3614));
    InMux I__714 (
            .O(N__3649),
            .I(N__3609));
    InMux I__713 (
            .O(N__3646),
            .I(N__3609));
    LocalMux I__712 (
            .O(N__3641),
            .I(ctrl_tap_fsm_state_2));
    LocalMux I__711 (
            .O(N__3636),
            .I(ctrl_tap_fsm_state_2));
    LocalMux I__710 (
            .O(N__3627),
            .I(ctrl_tap_fsm_state_2));
    Odrv4 I__709 (
            .O(N__3624),
            .I(ctrl_tap_fsm_state_2));
    LocalMux I__708 (
            .O(N__3619),
            .I(ctrl_tap_fsm_state_2));
    Odrv4 I__707 (
            .O(N__3614),
            .I(ctrl_tap_fsm_state_2));
    LocalMux I__706 (
            .O(N__3609),
            .I(ctrl_tap_fsm_state_2));
    CEMux I__705 (
            .O(N__3594),
            .I(N__3591));
    LocalMux I__704 (
            .O(N__3591),
            .I(N__3587));
    CEMux I__703 (
            .O(N__3590),
            .I(N__3584));
    Span4Mux_s1_v I__702 (
            .O(N__3587),
            .I(N__3579));
    LocalMux I__701 (
            .O(N__3584),
            .I(N__3579));
    Span4Mux_h I__700 (
            .O(N__3579),
            .I(N__3576));
    Odrv4 I__699 (
            .O(N__3576),
            .I(n1067));
    CascadeMux I__698 (
            .O(N__3573),
            .I(N__3570));
    InMux I__697 (
            .O(N__3570),
            .I(N__3567));
    LocalMux I__696 (
            .O(N__3567),
            .I(N__3563));
    InMux I__695 (
            .O(N__3566),
            .I(N__3560));
    Odrv12 I__694 (
            .O(N__3563),
            .I(ctrl_idcodeArea_shifter_22));
    LocalMux I__693 (
            .O(N__3560),
            .I(ctrl_idcodeArea_shifter_22));
    InMux I__692 (
            .O(N__3555),
            .I(N__3549));
    InMux I__691 (
            .O(N__3554),
            .I(N__3549));
    LocalMux I__690 (
            .O(N__3549),
            .I(ctrl_idcodeArea_shifter_21));
    IoInMux I__689 (
            .O(N__3546),
            .I(N__3543));
    LocalMux I__688 (
            .O(N__3543),
            .I(N__3540));
    Span4Mux_s1_h I__687 (
            .O(N__3540),
            .I(N__3536));
    InMux I__686 (
            .O(N__3539),
            .I(N__3533));
    Sp12to4 I__685 (
            .O(N__3536),
            .I(N__3529));
    LocalMux I__684 (
            .O(N__3533),
            .I(N__3526));
    InMux I__683 (
            .O(N__3532),
            .I(N__3523));
    Span12Mux_v I__682 (
            .O(N__3529),
            .I(N__3520));
    Span4Mux_v I__681 (
            .O(N__3526),
            .I(N__3515));
    LocalMux I__680 (
            .O(N__3523),
            .I(N__3515));
    Odrv12 I__679 (
            .O(N__3520),
            .I(io_leds_c_0));
    Odrv4 I__678 (
            .O(N__3515),
            .I(io_leds_c_0));
    InMux I__677 (
            .O(N__3510),
            .I(N__3506));
    InMux I__676 (
            .O(N__3509),
            .I(N__3503));
    LocalMux I__675 (
            .O(N__3506),
            .I(N__3500));
    LocalMux I__674 (
            .O(N__3503),
            .I(N__3497));
    Span4Mux_s3_v I__673 (
            .O(N__3500),
            .I(N__3494));
    Span4Mux_s3_h I__672 (
            .O(N__3497),
            .I(N__3491));
    Odrv4 I__671 (
            .O(N__3494),
            .I(ctrl_ledsArea_shifter_0));
    Odrv4 I__670 (
            .O(N__3491),
            .I(ctrl_ledsArea_shifter_0));
    SRMux I__669 (
            .O(N__3486),
            .I(N__3482));
    SRMux I__668 (
            .O(N__3485),
            .I(N__3479));
    LocalMux I__667 (
            .O(N__3482),
            .I(N__3475));
    LocalMux I__666 (
            .O(N__3479),
            .I(N__3472));
    SRMux I__665 (
            .O(N__3478),
            .I(N__3469));
    Span4Mux_v I__664 (
            .O(N__3475),
            .I(N__3464));
    Span4Mux_h I__663 (
            .O(N__3472),
            .I(N__3464));
    LocalMux I__662 (
            .O(N__3469),
            .I(N__3460));
    Span4Mux_v I__661 (
            .O(N__3464),
            .I(N__3457));
    SRMux I__660 (
            .O(N__3463),
            .I(N__3454));
    Span4Mux_v I__659 (
            .O(N__3460),
            .I(N__3451));
    Span4Mux_v I__658 (
            .O(N__3457),
            .I(N__3448));
    LocalMux I__657 (
            .O(N__3454),
            .I(N__3445));
    Span4Mux_v I__656 (
            .O(N__3451),
            .I(N__3442));
    Odrv4 I__655 (
            .O(N__3448),
            .I(global_reset_c));
    Odrv12 I__654 (
            .O(N__3445),
            .I(global_reset_c));
    Odrv4 I__653 (
            .O(N__3442),
            .I(global_reset_c));
    InMux I__652 (
            .O(N__3435),
            .I(N__3432));
    LocalMux I__651 (
            .O(N__3432),
            .I(N__3425));
    InMux I__650 (
            .O(N__3431),
            .I(N__3422));
    InMux I__649 (
            .O(N__3430),
            .I(N__3417));
    InMux I__648 (
            .O(N__3429),
            .I(N__3417));
    InMux I__647 (
            .O(N__3428),
            .I(N__3414));
    Odrv4 I__646 (
            .O(N__3425),
            .I(ctrl_tap_instruction_1));
    LocalMux I__645 (
            .O(N__3422),
            .I(ctrl_tap_instruction_1));
    LocalMux I__644 (
            .O(N__3417),
            .I(ctrl_tap_instruction_1));
    LocalMux I__643 (
            .O(N__3414),
            .I(ctrl_tap_instruction_1));
    CascadeMux I__642 (
            .O(N__3405),
            .I(N__3401));
    InMux I__641 (
            .O(N__3404),
            .I(N__3398));
    InMux I__640 (
            .O(N__3401),
            .I(N__3393));
    LocalMux I__639 (
            .O(N__3398),
            .I(N__3390));
    InMux I__638 (
            .O(N__3397),
            .I(N__3387));
    InMux I__637 (
            .O(N__3396),
            .I(N__3384));
    LocalMux I__636 (
            .O(N__3393),
            .I(ctrl_tap_instruction_2));
    Odrv4 I__635 (
            .O(N__3390),
            .I(ctrl_tap_instruction_2));
    LocalMux I__634 (
            .O(N__3387),
            .I(ctrl_tap_instruction_2));
    LocalMux I__633 (
            .O(N__3384),
            .I(ctrl_tap_instruction_2));
    InMux I__632 (
            .O(N__3375),
            .I(N__3372));
    LocalMux I__631 (
            .O(N__3372),
            .I(N__3368));
    InMux I__630 (
            .O(N__3371),
            .I(N__3365));
    Odrv12 I__629 (
            .O(N__3368),
            .I(ctrl_tap_instructionShift_2));
    LocalMux I__628 (
            .O(N__3365),
            .I(ctrl_tap_instructionShift_2));
    InMux I__627 (
            .O(N__3360),
            .I(N__3356));
    InMux I__626 (
            .O(N__3359),
            .I(N__3353));
    LocalMux I__625 (
            .O(N__3356),
            .I(N__3347));
    LocalMux I__624 (
            .O(N__3353),
            .I(N__3347));
    InMux I__623 (
            .O(N__3352),
            .I(N__3344));
    Odrv4 I__622 (
            .O(N__3347),
            .I(ctrl_tap_instruction_4));
    LocalMux I__621 (
            .O(N__3344),
            .I(ctrl_tap_instruction_4));
    InMux I__620 (
            .O(N__3339),
            .I(N__3336));
    LocalMux I__619 (
            .O(N__3336),
            .I(N__3331));
    InMux I__618 (
            .O(N__3335),
            .I(N__3326));
    InMux I__617 (
            .O(N__3334),
            .I(N__3326));
    Odrv12 I__616 (
            .O(N__3331),
            .I(ctrl_tap_instruction_5));
    LocalMux I__615 (
            .O(N__3326),
            .I(ctrl_tap_instruction_5));
    CascadeMux I__614 (
            .O(N__3321),
            .I(N__3318));
    InMux I__613 (
            .O(N__3318),
            .I(N__3315));
    LocalMux I__612 (
            .O(N__3315),
            .I(N__3312));
    Span4Mux_s2_h I__611 (
            .O(N__3312),
            .I(N__3308));
    InMux I__610 (
            .O(N__3311),
            .I(N__3305));
    Odrv4 I__609 (
            .O(N__3308),
            .I(ctrl_tap_instructionShift_5));
    LocalMux I__608 (
            .O(N__3305),
            .I(ctrl_tap_instructionShift_5));
    CascadeMux I__607 (
            .O(N__3300),
            .I(N__3296));
    InMux I__606 (
            .O(N__3299),
            .I(N__3293));
    InMux I__605 (
            .O(N__3296),
            .I(N__3288));
    LocalMux I__604 (
            .O(N__3293),
            .I(N__3285));
    InMux I__603 (
            .O(N__3292),
            .I(N__3280));
    InMux I__602 (
            .O(N__3291),
            .I(N__3280));
    LocalMux I__601 (
            .O(N__3288),
            .I(ctrl_tap_instruction_7));
    Odrv4 I__600 (
            .O(N__3285),
            .I(ctrl_tap_instruction_7));
    LocalMux I__599 (
            .O(N__3280),
            .I(ctrl_tap_instruction_7));
    CascadeMux I__598 (
            .O(N__3273),
            .I(N__3270));
    InMux I__597 (
            .O(N__3270),
            .I(N__3267));
    LocalMux I__596 (
            .O(N__3267),
            .I(N__3264));
    Span4Mux_s2_h I__595 (
            .O(N__3264),
            .I(N__3260));
    InMux I__594 (
            .O(N__3263),
            .I(N__3257));
    Odrv4 I__593 (
            .O(N__3260),
            .I(ctrl_tap_instructionShift_4));
    LocalMux I__592 (
            .O(N__3257),
            .I(ctrl_tap_instructionShift_4));
    InMux I__591 (
            .O(N__3252),
            .I(N__3248));
    CascadeMux I__590 (
            .O(N__3251),
            .I(N__3244));
    LocalMux I__589 (
            .O(N__3248),
            .I(N__3240));
    InMux I__588 (
            .O(N__3247),
            .I(N__3237));
    InMux I__587 (
            .O(N__3244),
            .I(N__3232));
    InMux I__586 (
            .O(N__3243),
            .I(N__3232));
    Odrv4 I__585 (
            .O(N__3240),
            .I(ctrl_tap_instruction_3));
    LocalMux I__584 (
            .O(N__3237),
            .I(ctrl_tap_instruction_3));
    LocalMux I__583 (
            .O(N__3232),
            .I(ctrl_tap_instruction_3));
    CascadeMux I__582 (
            .O(N__3225),
            .I(N__3222));
    InMux I__581 (
            .O(N__3222),
            .I(N__3219));
    LocalMux I__580 (
            .O(N__3219),
            .I(N__3215));
    InMux I__579 (
            .O(N__3218),
            .I(N__3212));
    Odrv4 I__578 (
            .O(N__3215),
            .I(ctrl_tap_instructionShift_3));
    LocalMux I__577 (
            .O(N__3212),
            .I(ctrl_tap_instructionShift_3));
    InMux I__576 (
            .O(N__3207),
            .I(N__3204));
    LocalMux I__575 (
            .O(N__3204),
            .I(N__3200));
    InMux I__574 (
            .O(N__3203),
            .I(N__3197));
    Odrv4 I__573 (
            .O(N__3200),
            .I(ctrl_tap_instructionShift_7));
    LocalMux I__572 (
            .O(N__3197),
            .I(ctrl_tap_instructionShift_7));
    InMux I__571 (
            .O(N__3192),
            .I(N__3189));
    LocalMux I__570 (
            .O(N__3189),
            .I(N__3183));
    InMux I__569 (
            .O(N__3188),
            .I(N__3176));
    InMux I__568 (
            .O(N__3187),
            .I(N__3176));
    InMux I__567 (
            .O(N__3186),
            .I(N__3176));
    Odrv12 I__566 (
            .O(N__3183),
            .I(ctrl_tap_instruction_6));
    LocalMux I__565 (
            .O(N__3176),
            .I(ctrl_tap_instruction_6));
    CascadeMux I__564 (
            .O(N__3171),
            .I(N__3168));
    InMux I__563 (
            .O(N__3168),
            .I(N__3165));
    LocalMux I__562 (
            .O(N__3165),
            .I(N__3161));
    InMux I__561 (
            .O(N__3164),
            .I(N__3158));
    Odrv4 I__560 (
            .O(N__3161),
            .I(ctrl_tap_instructionShift_6));
    LocalMux I__559 (
            .O(N__3158),
            .I(ctrl_tap_instructionShift_6));
    CascadeMux I__558 (
            .O(N__3153),
            .I(N__3150));
    InMux I__557 (
            .O(N__3150),
            .I(N__3147));
    LocalMux I__556 (
            .O(N__3147),
            .I(N__3143));
    InMux I__555 (
            .O(N__3146),
            .I(N__3140));
    Odrv12 I__554 (
            .O(N__3143),
            .I(ctrl_tap_instructionShift_1));
    LocalMux I__553 (
            .O(N__3140),
            .I(ctrl_tap_instructionShift_1));
    InMux I__552 (
            .O(N__3135),
            .I(N__3132));
    LocalMux I__551 (
            .O(N__3132),
            .I(N__3129));
    Span4Mux_h I__550 (
            .O(N__3129),
            .I(N__3122));
    InMux I__549 (
            .O(N__3128),
            .I(N__3119));
    InMux I__548 (
            .O(N__3127),
            .I(N__3116));
    InMux I__547 (
            .O(N__3126),
            .I(N__3113));
    InMux I__546 (
            .O(N__3125),
            .I(N__3110));
    Odrv4 I__545 (
            .O(N__3122),
            .I(ctrl_tap_instruction_0));
    LocalMux I__544 (
            .O(N__3119),
            .I(ctrl_tap_instruction_0));
    LocalMux I__543 (
            .O(N__3116),
            .I(ctrl_tap_instruction_0));
    LocalMux I__542 (
            .O(N__3113),
            .I(ctrl_tap_instruction_0));
    LocalMux I__541 (
            .O(N__3110),
            .I(ctrl_tap_instruction_0));
    CascadeMux I__540 (
            .O(N__3099),
            .I(N__3096));
    InMux I__539 (
            .O(N__3096),
            .I(N__3093));
    LocalMux I__538 (
            .O(N__3093),
            .I(N__3089));
    InMux I__537 (
            .O(N__3092),
            .I(N__3086));
    Span4Mux_s1_v I__536 (
            .O(N__3089),
            .I(N__3081));
    LocalMux I__535 (
            .O(N__3086),
            .I(N__3081));
    Odrv4 I__534 (
            .O(N__3081),
            .I(ctrl_tap_instructionShift_0));
    CascadeMux I__533 (
            .O(N__3078),
            .I(N__3075));
    InMux I__532 (
            .O(N__3075),
            .I(N__3069));
    InMux I__531 (
            .O(N__3074),
            .I(N__3069));
    LocalMux I__530 (
            .O(N__3069),
            .I(ctrl_idcodeArea_shifter_11));
    InMux I__529 (
            .O(N__3066),
            .I(N__3060));
    InMux I__528 (
            .O(N__3065),
            .I(N__3060));
    LocalMux I__527 (
            .O(N__3060),
            .I(ctrl_idcodeArea_shifter_10));
    InMux I__526 (
            .O(N__3057),
            .I(N__3053));
    InMux I__525 (
            .O(N__3056),
            .I(N__3050));
    LocalMux I__524 (
            .O(N__3053),
            .I(myClockArea_timeout_counter_value_4));
    LocalMux I__523 (
            .O(N__3050),
            .I(myClockArea_timeout_counter_value_4));
    InMux I__522 (
            .O(N__3045),
            .I(N__3041));
    InMux I__521 (
            .O(N__3044),
            .I(N__3038));
    LocalMux I__520 (
            .O(N__3041),
            .I(myClockArea_timeout_counter_value_6));
    LocalMux I__519 (
            .O(N__3038),
            .I(myClockArea_timeout_counter_value_6));
    CascadeMux I__518 (
            .O(N__3033),
            .I(N__3029));
    InMux I__517 (
            .O(N__3032),
            .I(N__3026));
    InMux I__516 (
            .O(N__3029),
            .I(N__3023));
    LocalMux I__515 (
            .O(N__3026),
            .I(myClockArea_timeout_counter_value_22));
    LocalMux I__514 (
            .O(N__3023),
            .I(myClockArea_timeout_counter_value_22));
    InMux I__513 (
            .O(N__3018),
            .I(N__3014));
    InMux I__512 (
            .O(N__3017),
            .I(N__3011));
    LocalMux I__511 (
            .O(N__3014),
            .I(myClockArea_timeout_counter_value_16));
    LocalMux I__510 (
            .O(N__3011),
            .I(myClockArea_timeout_counter_value_16));
    InMux I__509 (
            .O(N__3006),
            .I(N__3002));
    InMux I__508 (
            .O(N__3005),
            .I(N__2999));
    LocalMux I__507 (
            .O(N__3002),
            .I(myClockArea_timeout_counter_value_17));
    LocalMux I__506 (
            .O(N__2999),
            .I(myClockArea_timeout_counter_value_17));
    InMux I__505 (
            .O(N__2994),
            .I(N__2990));
    InMux I__504 (
            .O(N__2993),
            .I(N__2987));
    LocalMux I__503 (
            .O(N__2990),
            .I(myClockArea_timeout_counter_value_8));
    LocalMux I__502 (
            .O(N__2987),
            .I(myClockArea_timeout_counter_value_8));
    CascadeMux I__501 (
            .O(N__2982),
            .I(N__2978));
    InMux I__500 (
            .O(N__2981),
            .I(N__2975));
    InMux I__499 (
            .O(N__2978),
            .I(N__2972));
    LocalMux I__498 (
            .O(N__2975),
            .I(myClockArea_timeout_counter_value_10));
    LocalMux I__497 (
            .O(N__2972),
            .I(myClockArea_timeout_counter_value_10));
    InMux I__496 (
            .O(N__2967),
            .I(N__2963));
    InMux I__495 (
            .O(N__2966),
            .I(N__2960));
    LocalMux I__494 (
            .O(N__2963),
            .I(myClockArea_timeout_counter_value_2));
    LocalMux I__493 (
            .O(N__2960),
            .I(myClockArea_timeout_counter_value_2));
    InMux I__492 (
            .O(N__2955),
            .I(N__2952));
    LocalMux I__491 (
            .O(N__2952),
            .I(n2176));
    CascadeMux I__490 (
            .O(N__2949),
            .I(n2160_cascade_));
    InMux I__489 (
            .O(N__2946),
            .I(N__2943));
    LocalMux I__488 (
            .O(N__2943),
            .I(n2164));
    InMux I__487 (
            .O(N__2940),
            .I(N__2936));
    InMux I__486 (
            .O(N__2939),
            .I(N__2933));
    LocalMux I__485 (
            .O(N__2936),
            .I(myClockArea_timeout_counter_value_13));
    LocalMux I__484 (
            .O(N__2933),
            .I(myClockArea_timeout_counter_value_13));
    InMux I__483 (
            .O(N__2928),
            .I(N__2925));
    LocalMux I__482 (
            .O(N__2925),
            .I(n11));
    CascadeMux I__481 (
            .O(N__2922),
            .I(n2182_cascade_));
    InMux I__480 (
            .O(N__2919),
            .I(N__2916));
    LocalMux I__479 (
            .O(N__2916),
            .I(n13));
    CascadeMux I__478 (
            .O(N__2913),
            .I(n2113_cascade_));
    InMux I__477 (
            .O(N__2910),
            .I(N__2890));
    InMux I__476 (
            .O(N__2909),
            .I(N__2890));
    InMux I__475 (
            .O(N__2908),
            .I(N__2890));
    InMux I__474 (
            .O(N__2907),
            .I(N__2890));
    InMux I__473 (
            .O(N__2906),
            .I(N__2881));
    InMux I__472 (
            .O(N__2905),
            .I(N__2881));
    InMux I__471 (
            .O(N__2904),
            .I(N__2881));
    InMux I__470 (
            .O(N__2903),
            .I(N__2881));
    InMux I__469 (
            .O(N__2902),
            .I(N__2861));
    InMux I__468 (
            .O(N__2901),
            .I(N__2861));
    InMux I__467 (
            .O(N__2900),
            .I(N__2861));
    InMux I__466 (
            .O(N__2899),
            .I(N__2861));
    LocalMux I__465 (
            .O(N__2890),
            .I(N__2858));
    LocalMux I__464 (
            .O(N__2881),
            .I(N__2855));
    InMux I__463 (
            .O(N__2880),
            .I(N__2846));
    InMux I__462 (
            .O(N__2879),
            .I(N__2846));
    InMux I__461 (
            .O(N__2878),
            .I(N__2846));
    InMux I__460 (
            .O(N__2877),
            .I(N__2846));
    InMux I__459 (
            .O(N__2876),
            .I(N__2839));
    InMux I__458 (
            .O(N__2875),
            .I(N__2839));
    InMux I__457 (
            .O(N__2874),
            .I(N__2839));
    InMux I__456 (
            .O(N__2873),
            .I(N__2830));
    InMux I__455 (
            .O(N__2872),
            .I(N__2830));
    InMux I__454 (
            .O(N__2871),
            .I(N__2830));
    InMux I__453 (
            .O(N__2870),
            .I(N__2830));
    LocalMux I__452 (
            .O(N__2861),
            .I(n1771));
    Odrv4 I__451 (
            .O(N__2858),
            .I(n1771));
    Odrv4 I__450 (
            .O(N__2855),
            .I(n1771));
    LocalMux I__449 (
            .O(N__2846),
            .I(n1771));
    LocalMux I__448 (
            .O(N__2839),
            .I(n1771));
    LocalMux I__447 (
            .O(N__2830),
            .I(n1771));
    InMux I__446 (
            .O(N__2817),
            .I(N__2813));
    InMux I__445 (
            .O(N__2816),
            .I(N__2810));
    LocalMux I__444 (
            .O(N__2813),
            .I(myClockArea_timeout_counter_value_19));
    LocalMux I__443 (
            .O(N__2810),
            .I(myClockArea_timeout_counter_value_19));
    InMux I__442 (
            .O(N__2805),
            .I(N__2801));
    InMux I__441 (
            .O(N__2804),
            .I(N__2798));
    LocalMux I__440 (
            .O(N__2801),
            .I(myClockArea_timeout_counter_value_15));
    LocalMux I__439 (
            .O(N__2798),
            .I(myClockArea_timeout_counter_value_15));
    CascadeMux I__438 (
            .O(N__2793),
            .I(N__2789));
    InMux I__437 (
            .O(N__2792),
            .I(N__2786));
    InMux I__436 (
            .O(N__2789),
            .I(N__2783));
    LocalMux I__435 (
            .O(N__2786),
            .I(myClockArea_timeout_counter_value_20));
    LocalMux I__434 (
            .O(N__2783),
            .I(myClockArea_timeout_counter_value_20));
    InMux I__433 (
            .O(N__2778),
            .I(N__2774));
    InMux I__432 (
            .O(N__2777),
            .I(N__2771));
    LocalMux I__431 (
            .O(N__2774),
            .I(myClockArea_timeout_counter_value_11));
    LocalMux I__430 (
            .O(N__2771),
            .I(myClockArea_timeout_counter_value_11));
    InMux I__429 (
            .O(N__2766),
            .I(N__2763));
    LocalMux I__428 (
            .O(N__2763),
            .I(n2162));
    InMux I__427 (
            .O(N__2760),
            .I(N__2757));
    LocalMux I__426 (
            .O(N__2757),
            .I(n2113));
    InMux I__425 (
            .O(N__2754),
            .I(N__2737));
    InMux I__424 (
            .O(N__2753),
            .I(N__2737));
    InMux I__423 (
            .O(N__2752),
            .I(N__2737));
    InMux I__422 (
            .O(N__2751),
            .I(N__2737));
    InMux I__421 (
            .O(N__2750),
            .I(N__2737));
    InMux I__420 (
            .O(N__2749),
            .I(N__2734));
    InMux I__419 (
            .O(N__2748),
            .I(N__2731));
    LocalMux I__418 (
            .O(N__2737),
            .I(n12_adj_3));
    LocalMux I__417 (
            .O(N__2734),
            .I(n12_adj_3));
    LocalMux I__416 (
            .O(N__2731),
            .I(n12_adj_3));
    InMux I__415 (
            .O(N__2724),
            .I(N__2712));
    InMux I__414 (
            .O(N__2723),
            .I(N__2712));
    InMux I__413 (
            .O(N__2722),
            .I(N__2712));
    InMux I__412 (
            .O(N__2721),
            .I(N__2712));
    LocalMux I__411 (
            .O(N__2712),
            .I(n1769));
    InMux I__410 (
            .O(N__2709),
            .I(N__2706));
    LocalMux I__409 (
            .O(N__2706),
            .I(n1864));
    InMux I__408 (
            .O(N__2703),
            .I(N__2699));
    InMux I__407 (
            .O(N__2702),
            .I(N__2696));
    LocalMux I__406 (
            .O(N__2699),
            .I(myClockArea_timeout_counter_value_3));
    LocalMux I__405 (
            .O(N__2696),
            .I(myClockArea_timeout_counter_value_3));
    InMux I__404 (
            .O(N__2691),
            .I(N__2687));
    InMux I__403 (
            .O(N__2690),
            .I(N__2684));
    LocalMux I__402 (
            .O(N__2687),
            .I(myClockArea_timeout_counter_value_1));
    LocalMux I__401 (
            .O(N__2684),
            .I(myClockArea_timeout_counter_value_1));
    CascadeMux I__400 (
            .O(N__2679),
            .I(N__2675));
    InMux I__399 (
            .O(N__2678),
            .I(N__2672));
    InMux I__398 (
            .O(N__2675),
            .I(N__2669));
    LocalMux I__397 (
            .O(N__2672),
            .I(myClockArea_timeout_counter_value_5));
    LocalMux I__396 (
            .O(N__2669),
            .I(myClockArea_timeout_counter_value_5));
    InMux I__395 (
            .O(N__2664),
            .I(N__2660));
    InMux I__394 (
            .O(N__2663),
            .I(N__2657));
    LocalMux I__393 (
            .O(N__2660),
            .I(myClockArea_timeout_counter_value_0));
    LocalMux I__392 (
            .O(N__2657),
            .I(myClockArea_timeout_counter_value_0));
    InMux I__391 (
            .O(N__2652),
            .I(N__2648));
    InMux I__390 (
            .O(N__2651),
            .I(N__2645));
    LocalMux I__389 (
            .O(N__2648),
            .I(myClockArea_timeout_counter_value_9));
    LocalMux I__388 (
            .O(N__2645),
            .I(myClockArea_timeout_counter_value_9));
    InMux I__387 (
            .O(N__2640),
            .I(N__2636));
    InMux I__386 (
            .O(N__2639),
            .I(N__2633));
    LocalMux I__385 (
            .O(N__2636),
            .I(N__2630));
    LocalMux I__384 (
            .O(N__2633),
            .I(myClockArea_timeout_counter_value_18));
    Odrv4 I__383 (
            .O(N__2630),
            .I(myClockArea_timeout_counter_value_18));
    CascadeMux I__382 (
            .O(N__2625),
            .I(N__2621));
    InMux I__381 (
            .O(N__2624),
            .I(N__2618));
    InMux I__380 (
            .O(N__2621),
            .I(N__2615));
    LocalMux I__379 (
            .O(N__2618),
            .I(myClockArea_timeout_counter_value_12));
    LocalMux I__378 (
            .O(N__2615),
            .I(myClockArea_timeout_counter_value_12));
    InMux I__377 (
            .O(N__2610),
            .I(N__2606));
    InMux I__376 (
            .O(N__2609),
            .I(N__2603));
    LocalMux I__375 (
            .O(N__2606),
            .I(myClockArea_timeout_counter_value_14));
    LocalMux I__374 (
            .O(N__2603),
            .I(myClockArea_timeout_counter_value_14));
    CascadeMux I__373 (
            .O(N__2598),
            .I(N__2594));
    InMux I__372 (
            .O(N__2597),
            .I(N__2591));
    InMux I__371 (
            .O(N__2594),
            .I(N__2588));
    LocalMux I__370 (
            .O(N__2591),
            .I(ctrl_idcodeArea_shifter_9));
    LocalMux I__369 (
            .O(N__2588),
            .I(ctrl_idcodeArea_shifter_9));
    InMux I__368 (
            .O(N__2583),
            .I(N__2579));
    InMux I__367 (
            .O(N__2582),
            .I(N__2576));
    LocalMux I__366 (
            .O(N__2579),
            .I(myClockArea_timeout_counter_value_7));
    LocalMux I__365 (
            .O(N__2576),
            .I(myClockArea_timeout_counter_value_7));
    InMux I__364 (
            .O(N__2571),
            .I(N__2567));
    InMux I__363 (
            .O(N__2570),
            .I(N__2564));
    LocalMux I__362 (
            .O(N__2567),
            .I(N__2561));
    LocalMux I__361 (
            .O(N__2564),
            .I(myClockArea_timeout_counter_value_21));
    Odrv4 I__360 (
            .O(N__2561),
            .I(myClockArea_timeout_counter_value_21));
    CascadeMux I__359 (
            .O(N__2556),
            .I(N__2552));
    InMux I__358 (
            .O(N__2555),
            .I(N__2549));
    InMux I__357 (
            .O(N__2552),
            .I(N__2546));
    LocalMux I__356 (
            .O(N__2549),
            .I(ctrl_idcodeArea_shifter_5));
    LocalMux I__355 (
            .O(N__2546),
            .I(ctrl_idcodeArea_shifter_5));
    CascadeMux I__354 (
            .O(N__2541),
            .I(N__2537));
    InMux I__353 (
            .O(N__2540),
            .I(N__2532));
    InMux I__352 (
            .O(N__2537),
            .I(N__2532));
    LocalMux I__351 (
            .O(N__2532),
            .I(ctrl_idcodeArea_shifter_7));
    CascadeMux I__350 (
            .O(N__2529),
            .I(N__2525));
    InMux I__349 (
            .O(N__2528),
            .I(N__2522));
    InMux I__348 (
            .O(N__2525),
            .I(N__2519));
    LocalMux I__347 (
            .O(N__2522),
            .I(ctrl_idcodeArea_shifter_6));
    LocalMux I__346 (
            .O(N__2519),
            .I(ctrl_idcodeArea_shifter_6));
    InMux I__345 (
            .O(N__2514),
            .I(N__2497));
    InMux I__344 (
            .O(N__2513),
            .I(N__2497));
    InMux I__343 (
            .O(N__2512),
            .I(N__2497));
    InMux I__342 (
            .O(N__2511),
            .I(N__2497));
    InMux I__341 (
            .O(N__2510),
            .I(N__2497));
    InMux I__340 (
            .O(N__2509),
            .I(N__2492));
    InMux I__339 (
            .O(N__2508),
            .I(N__2492));
    LocalMux I__338 (
            .O(N__2497),
            .I(n2045));
    LocalMux I__337 (
            .O(N__2492),
            .I(n2045));
    CascadeMux I__336 (
            .O(N__2487),
            .I(N__2483));
    InMux I__335 (
            .O(N__2486),
            .I(N__2480));
    InMux I__334 (
            .O(N__2483),
            .I(N__2477));
    LocalMux I__333 (
            .O(N__2480),
            .I(ctrl_idcodeArea_shifter_8));
    LocalMux I__332 (
            .O(N__2477),
            .I(ctrl_idcodeArea_shifter_8));
    InMux I__331 (
            .O(N__2472),
            .I(N__2469));
    LocalMux I__330 (
            .O(N__2469),
            .I(n2140));
    CascadeMux I__329 (
            .O(N__2466),
            .I(n9_cascade_));
    InMux I__328 (
            .O(N__2463),
            .I(N__2460));
    LocalMux I__327 (
            .O(N__2460),
            .I(n2191));
    InMux I__326 (
            .O(N__2457),
            .I(N__2453));
    InMux I__325 (
            .O(N__2456),
            .I(N__2450));
    LocalMux I__324 (
            .O(N__2453),
            .I(ctrl_idcodeArea_shifter_25));
    LocalMux I__323 (
            .O(N__2450),
            .I(ctrl_idcodeArea_shifter_25));
    InMux I__322 (
            .O(N__2445),
            .I(N__2442));
    LocalMux I__321 (
            .O(N__2442),
            .I(n6));
    InMux I__320 (
            .O(N__2439),
            .I(N__2435));
    InMux I__319 (
            .O(N__2438),
            .I(N__2432));
    LocalMux I__318 (
            .O(N__2435),
            .I(n1293));
    LocalMux I__317 (
            .O(N__2432),
            .I(n1293));
    CascadeMux I__316 (
            .O(N__2427),
            .I(n1582_cascade_));
    InMux I__315 (
            .O(N__2424),
            .I(N__2420));
    InMux I__314 (
            .O(N__2423),
            .I(N__2417));
    LocalMux I__313 (
            .O(N__2420),
            .I(n2119));
    LocalMux I__312 (
            .O(N__2417),
            .I(n2119));
    InMux I__311 (
            .O(N__2412),
            .I(N__2406));
    InMux I__310 (
            .O(N__2411),
            .I(N__2406));
    LocalMux I__309 (
            .O(N__2406),
            .I(ctrl_idcodeArea_shifter_24));
    CascadeMux I__308 (
            .O(N__2403),
            .I(n2178_cascade_));
    InMux I__307 (
            .O(N__2400),
            .I(N__2394));
    InMux I__306 (
            .O(N__2399),
            .I(N__2394));
    LocalMux I__305 (
            .O(N__2394),
            .I(ctrl_idcodeArea_shifter_23));
    CascadeMux I__304 (
            .O(N__2391),
            .I(n1313_cascade_));
    InMux I__303 (
            .O(N__2388),
            .I(N__2385));
    LocalMux I__302 (
            .O(N__2385),
            .I(ctrl_tap_tdoUnbufferd_N_224));
    CascadeMux I__301 (
            .O(N__2382),
            .I(N__2378));
    CascadeMux I__300 (
            .O(N__2381),
            .I(N__2375));
    InMux I__299 (
            .O(N__2378),
            .I(N__2372));
    InMux I__298 (
            .O(N__2375),
            .I(N__2369));
    LocalMux I__297 (
            .O(N__2372),
            .I(ctrl_idcodeArea_shifter_1));
    LocalMux I__296 (
            .O(N__2369),
            .I(ctrl_idcodeArea_shifter_1));
    InMux I__295 (
            .O(N__2364),
            .I(N__2360));
    InMux I__294 (
            .O(N__2363),
            .I(N__2357));
    LocalMux I__293 (
            .O(N__2360),
            .I(N__2354));
    LocalMux I__292 (
            .O(N__2357),
            .I(ctrl_idcodeArea_shifter_0));
    Odrv4 I__291 (
            .O(N__2354),
            .I(ctrl_idcodeArea_shifter_0));
    CascadeMux I__290 (
            .O(N__2349),
            .I(N__2345));
    InMux I__289 (
            .O(N__2348),
            .I(N__2342));
    InMux I__288 (
            .O(N__2345),
            .I(N__2339));
    LocalMux I__287 (
            .O(N__2342),
            .I(ctrl_idcodeArea_shifter_29));
    LocalMux I__286 (
            .O(N__2339),
            .I(ctrl_idcodeArea_shifter_29));
    CascadeMux I__285 (
            .O(N__2334),
            .I(N__2331));
    InMux I__284 (
            .O(N__2331),
            .I(N__2325));
    InMux I__283 (
            .O(N__2330),
            .I(N__2325));
    LocalMux I__282 (
            .O(N__2325),
            .I(ctrl_idcodeArea_shifter_28));
    CascadeMux I__281 (
            .O(N__2322),
            .I(N__2319));
    InMux I__280 (
            .O(N__2319),
            .I(N__2313));
    InMux I__279 (
            .O(N__2318),
            .I(N__2313));
    LocalMux I__278 (
            .O(N__2313),
            .I(ctrl_idcodeArea_shifter_27));
    CascadeMux I__277 (
            .O(N__2310),
            .I(N__2307));
    InMux I__276 (
            .O(N__2307),
            .I(N__2301));
    InMux I__275 (
            .O(N__2306),
            .I(N__2301));
    LocalMux I__274 (
            .O(N__2301),
            .I(ctrl_idcodeArea_shifter_26));
    InMux I__273 (
            .O(N__2298),
            .I(n2030));
    InMux I__272 (
            .O(N__2295),
            .I(N__2292));
    LocalMux I__271 (
            .O(N__2292),
            .I(n2116));
    CascadeMux I__270 (
            .O(N__2289),
            .I(n4_cascade_));
    CascadeMux I__269 (
            .O(N__2286),
            .I(ctrl_tap_tdoUnbufferd_N_223_cascade_));
    IoInMux I__268 (
            .O(N__2283),
            .I(N__2280));
    LocalMux I__267 (
            .O(N__2280),
            .I(N__2277));
    IoSpan4Mux I__266 (
            .O(N__2277),
            .I(N__2274));
    Odrv4 I__265 (
            .O(N__2274),
            .I(ctrl_tap_tdoUnbufferd));
    InMux I__264 (
            .O(N__2271),
            .I(N__2261));
    InMux I__263 (
            .O(N__2270),
            .I(N__2256));
    InMux I__262 (
            .O(N__2269),
            .I(N__2256));
    InMux I__261 (
            .O(N__2268),
            .I(N__2245));
    InMux I__260 (
            .O(N__2267),
            .I(N__2245));
    InMux I__259 (
            .O(N__2266),
            .I(N__2245));
    InMux I__258 (
            .O(N__2265),
            .I(N__2245));
    InMux I__257 (
            .O(N__2264),
            .I(N__2245));
    LocalMux I__256 (
            .O(N__2261),
            .I(n2146));
    LocalMux I__255 (
            .O(N__2256),
            .I(n2146));
    LocalMux I__254 (
            .O(N__2245),
            .I(n2146));
    InMux I__253 (
            .O(N__2238),
            .I(n2021));
    InMux I__252 (
            .O(N__2235),
            .I(n2022));
    InMux I__251 (
            .O(N__2232),
            .I(n2023));
    InMux I__250 (
            .O(N__2229),
            .I(bfn_1_8_0_));
    InMux I__249 (
            .O(N__2226),
            .I(n2025));
    InMux I__248 (
            .O(N__2223),
            .I(n2026));
    InMux I__247 (
            .O(N__2220),
            .I(n2027));
    InMux I__246 (
            .O(N__2217),
            .I(n2028));
    InMux I__245 (
            .O(N__2214),
            .I(n2029));
    InMux I__244 (
            .O(N__2211),
            .I(n2012));
    InMux I__243 (
            .O(N__2208),
            .I(n2013));
    InMux I__242 (
            .O(N__2205),
            .I(n2014));
    InMux I__241 (
            .O(N__2202),
            .I(n2015));
    InMux I__240 (
            .O(N__2199),
            .I(bfn_1_7_0_));
    InMux I__239 (
            .O(N__2196),
            .I(n2017));
    InMux I__238 (
            .O(N__2193),
            .I(n2018));
    InMux I__237 (
            .O(N__2190),
            .I(n2019));
    InMux I__236 (
            .O(N__2187),
            .I(n2020));
    InMux I__235 (
            .O(N__2184),
            .I(N__2181));
    LocalMux I__234 (
            .O(N__2181),
            .I(n1023));
    InMux I__233 (
            .O(N__2178),
            .I(N__2174));
    InMux I__232 (
            .O(N__2177),
            .I(N__2171));
    LocalMux I__231 (
            .O(N__2174),
            .I(n1027));
    LocalMux I__230 (
            .O(N__2171),
            .I(n1027));
    InMux I__229 (
            .O(N__2166),
            .I(N__2163));
    LocalMux I__228 (
            .O(N__2163),
            .I(n965));
    InMux I__227 (
            .O(N__2160),
            .I(N__2157));
    LocalMux I__226 (
            .O(N__2157),
            .I(n5));
    CascadeMux I__225 (
            .O(N__2154),
            .I(n5_cascade_));
    InMux I__224 (
            .O(N__2151),
            .I(N__2148));
    LocalMux I__223 (
            .O(N__2148),
            .I(n2201));
    InMux I__222 (
            .O(N__2145),
            .I(bfn_1_6_0_));
    InMux I__221 (
            .O(N__2142),
            .I(n2009));
    InMux I__220 (
            .O(N__2139),
            .I(n2010));
    InMux I__219 (
            .O(N__2136),
            .I(n2011));
    CascadeMux I__218 (
            .O(N__2133),
            .I(n2188_cascade_));
    CascadeMux I__217 (
            .O(N__2130),
            .I(n2235_cascade_));
    CascadeMux I__216 (
            .O(N__2127),
            .I(n2202_cascade_));
    CascadeMux I__215 (
            .O(N__2124),
            .I(N__2121));
    InMux I__214 (
            .O(N__2121),
            .I(N__2118));
    LocalMux I__213 (
            .O(N__2118),
            .I(N__2115));
    Odrv12 I__212 (
            .O(N__2115),
            .I(n2211));
    InMux I__211 (
            .O(N__2112),
            .I(N__2109));
    LocalMux I__210 (
            .O(N__2109),
            .I(n962));
    InMux I__209 (
            .O(N__2106),
            .I(N__2103));
    LocalMux I__208 (
            .O(N__2103),
            .I(n1025));
    CascadeMux I__207 (
            .O(N__2100),
            .I(n1025_cascade_));
    CascadeMux I__206 (
            .O(N__2097),
            .I(n960_cascade_));
    InMux I__205 (
            .O(N__2094),
            .I(N__2091));
    LocalMux I__204 (
            .O(N__2091),
            .I(n2194));
    CascadeMux I__203 (
            .O(N__2088),
            .I(N__2085));
    InMux I__202 (
            .O(N__2085),
            .I(N__2082));
    LocalMux I__201 (
            .O(N__2082),
            .I(n1828));
    CascadeMux I__200 (
            .O(N__2079),
            .I(n2045_cascade_));
    CascadeMux I__199 (
            .O(N__2076),
            .I(N__2072));
    InMux I__198 (
            .O(N__2075),
            .I(N__2067));
    InMux I__197 (
            .O(N__2072),
            .I(N__2067));
    LocalMux I__196 (
            .O(N__2067),
            .I(ctrl_idcodeArea_shifter_4));
    CascadeMux I__195 (
            .O(N__2064),
            .I(N__2060));
    InMux I__194 (
            .O(N__2063),
            .I(N__2057));
    InMux I__193 (
            .O(N__2060),
            .I(N__2054));
    LocalMux I__192 (
            .O(N__2057),
            .I(ctrl_idcodeArea_shifter_3));
    LocalMux I__191 (
            .O(N__2054),
            .I(ctrl_idcodeArea_shifter_3));
    InMux I__190 (
            .O(N__2049),
            .I(N__2043));
    InMux I__189 (
            .O(N__2048),
            .I(N__2043));
    LocalMux I__188 (
            .O(N__2043),
            .I(ctrl_idcodeArea_shifter_30));
    CascadeMux I__187 (
            .O(N__2040),
            .I(n1854_cascade_));
    CascadeMux I__186 (
            .O(N__2037),
            .I(n9_adj_2_cascade_));
    InMux I__185 (
            .O(N__2034),
            .I(N__2031));
    LocalMux I__184 (
            .O(N__2031),
            .I(n8));
    InMux I__183 (
            .O(N__2028),
            .I(N__2025));
    LocalMux I__182 (
            .O(N__2025),
            .I(n12));
    CascadeMux I__181 (
            .O(N__2022),
            .I(n2_cascade_));
    InMux I__180 (
            .O(N__2019),
            .I(N__2013));
    InMux I__179 (
            .O(N__2018),
            .I(N__2013));
    LocalMux I__178 (
            .O(N__2013),
            .I(ctrl_idcodeArea_shifter_2));
    CascadeMux I__177 (
            .O(N__2010),
            .I(n12_cascade_));
    InMux I__176 (
            .O(N__2007),
            .I(N__2004));
    LocalMux I__175 (
            .O(N__2004),
            .I(n1307));
    CascadeMux I__174 (
            .O(N__2001),
            .I(n2116_cascade_));
    IoInMux I__173 (
            .O(N__1998),
            .I(N__1995));
    LocalMux I__172 (
            .O(N__1995),
            .I(N__1992));
    Span4Mux_s3_h I__171 (
            .O(N__1992),
            .I(N__1989));
    Sp12to4 I__170 (
            .O(N__1989),
            .I(N__1986));
    Odrv12 I__169 (
            .O(N__1986),
            .I(io_jtag_tck_pad_gb_input));
    defparam IN_MUX_bfv_1_6_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_6_0_));
    defparam IN_MUX_bfv_1_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_7_0_ (
            .carryinitin(n2016),
            .carryinitout(bfn_1_7_0_));
    defparam IN_MUX_bfv_1_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_8_0_ (
            .carryinitin(n2024),
            .carryinitout(bfn_1_8_0_));
    ICE_GB io_jtag_tck_pad_gb (
            .USERSIGNALTOGLOBALBUFFER(N__1998),
            .GLOBALBUFFEROUTPUT(io_jtag_tck_c));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam i1_2_lut_adj_4_LC_1_1_0.C_ON=1'b0;
    defparam i1_2_lut_adj_4_LC_1_1_0.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_4_LC_1_1_0.LUT_INIT=16'b1110111011101110;
    LogicCell40 i1_2_lut_adj_4_LC_1_1_0 (
            .in0(N__3291),
            .in1(N__3186),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(n1307),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_tap_instruction_i1_LC_1_1_1.C_ON=1'b0;
    defparam ctrl_tap_instruction_i1_LC_1_1_1.SEQ_MODE=4'b1000;
    defparam ctrl_tap_instruction_i1_LC_1_1_1.LUT_INIT=16'b1011100000000000;
    LogicCell40 ctrl_tap_instruction_i1_LC_1_1_1 (
            .in0(N__3430),
            .in1(N__2269),
            .in2(N__3153),
            .in3(N__4921),
            .lcout(ctrl_tap_instruction_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4707),
            .ce(),
            .sr(_gnd_net_));
    defparam equal_312_i15_2_lut_LC_1_1_2.C_ON=1'b0;
    defparam equal_312_i15_2_lut_LC_1_1_2.SEQ_MODE=4'b0000;
    defparam equal_312_i15_2_lut_LC_1_1_2.LUT_INIT=16'b1111111111001100;
    LogicCell40 equal_312_i15_2_lut_LC_1_1_2 (
            .in0(_gnd_net_),
            .in1(N__3352),
            .in2(_gnd_net_),
            .in3(N__3334),
            .lcout(n12),
            .ltout(n12_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_6_LC_1_1_3.C_ON=1'b0;
    defparam i1_4_lut_adj_6_LC_1_1_3.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_6_LC_1_1_3.LUT_INIT=16'b1111111111111011;
    LogicCell40 i1_4_lut_adj_6_LC_1_1_3 (
            .in0(N__3243),
            .in1(N__3396),
            .in2(N__2010),
            .in3(N__2007),
            .lcout(n2116),
            .ltout(n2116_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_adj_5_LC_1_1_4.C_ON=1'b0;
    defparam i1_2_lut_3_lut_adj_5_LC_1_1_4.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_adj_5_LC_1_1_4.LUT_INIT=16'b1111001111111111;
    LogicCell40 i1_2_lut_3_lut_adj_5_LC_1_1_4 (
            .in0(_gnd_net_),
            .in1(N__3429),
            .in2(N__2001),
            .in3(N__3126),
            .lcout(n15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_2_lut_3_lut_LC_1_1_5.C_ON=1'b0;
    defparam i2_2_lut_3_lut_LC_1_1_5.SEQ_MODE=4'b0000;
    defparam i2_2_lut_3_lut_LC_1_1_5.LUT_INIT=16'b1111111111111010;
    LogicCell40 i2_2_lut_3_lut_LC_1_1_5 (
            .in0(N__3187),
            .in1(_gnd_net_),
            .in2(N__3251),
            .in3(N__3292),
            .lcout(n8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_tap_instruction_i6_LC_1_1_6.C_ON=1'b0;
    defparam ctrl_tap_instruction_i6_LC_1_1_6.SEQ_MODE=4'b1000;
    defparam ctrl_tap_instruction_i6_LC_1_1_6.LUT_INIT=16'b1010100000100000;
    LogicCell40 ctrl_tap_instruction_i6_LC_1_1_6 (
            .in0(N__4920),
            .in1(N__2271),
            .in2(N__3171),
            .in3(N__3188),
            .lcout(ctrl_tap_instruction_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4707),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_tap_instruction_i5_LC_1_1_7.C_ON=1'b0;
    defparam ctrl_tap_instruction_i5_LC_1_1_7.SEQ_MODE=4'b1000;
    defparam ctrl_tap_instruction_i5_LC_1_1_7.LUT_INIT=16'b1011100000000000;
    LogicCell40 ctrl_tap_instruction_i5_LC_1_1_7 (
            .in0(N__3335),
            .in1(N__2270),
            .in2(N__3321),
            .in3(N__4922),
            .lcout(ctrl_tap_instruction_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4707),
            .ce(),
            .sr(_gnd_net_));
    defparam i1047_2_lut_LC_1_2_0.C_ON=1'b0;
    defparam i1047_2_lut_LC_1_2_0.SEQ_MODE=4'b0000;
    defparam i1047_2_lut_LC_1_2_0.LUT_INIT=16'b1000100010001000;
    LogicCell40 i1047_2_lut_LC_1_2_0 (
            .in0(N__3431),
            .in1(N__3127),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(n1828),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i20_3_lut_3_lut_LC_1_2_1.C_ON=1'b0;
    defparam i20_3_lut_3_lut_LC_1_2_1.SEQ_MODE=4'b0000;
    defparam i20_3_lut_3_lut_LC_1_2_1.LUT_INIT=16'b0000010110101010;
    LogicCell40 i20_3_lut_3_lut_LC_1_2_1 (
            .in0(N__3870),
            .in1(_gnd_net_),
            .in2(N__4214),
            .in3(N__3683),
            .lcout(),
            .ltout(n9_adj_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1424_3_lut_LC_1_2_2.C_ON=1'b0;
    defparam i1424_3_lut_LC_1_2_2.SEQ_MODE=4'b0000;
    defparam i1424_3_lut_LC_1_2_2.LUT_INIT=16'b1100110000001100;
    LogicCell40 i1424_3_lut_LC_1_2_2 (
            .in0(_gnd_net_),
            .in1(N__3937),
            .in2(N__2037),
            .in3(N__4076),
            .lcout(n2211),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_idcodeArea_shifter_i2_LC_1_2_3.C_ON=1'b0;
    defparam ctrl_idcodeArea_shifter_i2_LC_1_2_3.SEQ_MODE=4'b1000;
    defparam ctrl_idcodeArea_shifter_i2_LC_1_2_3.LUT_INIT=16'b1010110000000000;
    LogicCell40 ctrl_idcodeArea_shifter_i2_LC_1_2_3 (
            .in0(N__2018),
            .in1(N__2063),
            .in2(N__5082),
            .in3(N__4866),
            .lcout(ctrl_idcodeArea_shifter_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4705),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_1_LC_1_2_4.C_ON=1'b0;
    defparam i1_2_lut_adj_1_LC_1_2_4.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_1_LC_1_2_4.LUT_INIT=16'b1100110000000000;
    LogicCell40 i1_2_lut_adj_1_LC_1_2_4 (
            .in0(_gnd_net_),
            .in1(N__4184),
            .in2(_gnd_net_),
            .in3(N__3869),
            .lcout(),
            .ltout(n2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i5_4_lut_LC_1_2_5.C_ON=1'b0;
    defparam i5_4_lut_LC_1_2_5.SEQ_MODE=4'b0000;
    defparam i5_4_lut_LC_1_2_5.LUT_INIT=16'b1110111111111111;
    LogicCell40 i5_4_lut_LC_1_2_5 (
            .in0(N__2034),
            .in1(N__2028),
            .in2(N__2022),
            .in3(N__3397),
            .lcout(n1293),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1343_2_lut_3_lut_LC_1_2_6.C_ON=1'b0;
    defparam i1343_2_lut_3_lut_LC_1_2_6.SEQ_MODE=4'b0000;
    defparam i1343_2_lut_3_lut_LC_1_2_6.LUT_INIT=16'b1111111111101110;
    LogicCell40 i1343_2_lut_3_lut_LC_1_2_6 (
            .in0(N__3684),
            .in1(N__4188),
            .in2(_gnd_net_),
            .in3(N__3871),
            .lcout(n2146),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_idcodeArea_shifter_i1_LC_1_2_7.C_ON=1'b0;
    defparam ctrl_idcodeArea_shifter_i1_LC_1_2_7.SEQ_MODE=4'b1000;
    defparam ctrl_idcodeArea_shifter_i1_LC_1_2_7.LUT_INIT=16'b1100000010001000;
    LogicCell40 ctrl_idcodeArea_shifter_i1_LC_1_2_7 (
            .in0(N__2019),
            .in1(N__4865),
            .in2(N__2381),
            .in3(N__5078),
            .lcout(ctrl_idcodeArea_shifter_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4705),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_idcodeArea_shifter_i4_LC_1_3_0.C_ON=1'b0;
    defparam ctrl_idcodeArea_shifter_i4_LC_1_3_0.SEQ_MODE=4'b1000;
    defparam ctrl_idcodeArea_shifter_i4_LC_1_3_0.LUT_INIT=16'b1100000010001000;
    LogicCell40 ctrl_idcodeArea_shifter_i4_LC_1_3_0 (
            .in0(N__2555),
            .in1(N__4859),
            .in2(N__2076),
            .in3(N__5048),
            .lcout(ctrl_idcodeArea_shifter_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4703),
            .ce(),
            .sr(_gnd_net_));
    defparam i3_4_lut_LC_1_3_1.C_ON=1'b0;
    defparam i3_4_lut_LC_1_3_1.SEQ_MODE=4'b0000;
    defparam i3_4_lut_LC_1_3_1.LUT_INIT=16'b1011111111111111;
    LogicCell40 i3_4_lut_LC_1_3_1 (
            .in0(N__2438),
            .in1(N__3659),
            .in2(N__2088),
            .in3(N__4052),
            .lcout(n2045),
            .ltout(n2045_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_ledsArea_store_i0_i7_LC_1_3_2.C_ON=1'b0;
    defparam ctrl_ledsArea_store_i0_i7_LC_1_3_2.SEQ_MODE=4'b1000;
    defparam ctrl_ledsArea_store_i0_i7_LC_1_3_2.LUT_INIT=16'b1111101000001010;
    LogicCell40 ctrl_ledsArea_store_i0_i7_LC_1_3_2 (
            .in0(N__4392),
            .in1(_gnd_net_),
            .in2(N__2079),
            .in3(N__4408),
            .lcout(io_leds_c_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4703),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_idcodeArea_shifter_i3_LC_1_3_3.C_ON=1'b0;
    defparam ctrl_idcodeArea_shifter_i3_LC_1_3_3.SEQ_MODE=4'b1000;
    defparam ctrl_idcodeArea_shifter_i3_LC_1_3_3.LUT_INIT=16'b1110010000000000;
    LogicCell40 ctrl_idcodeArea_shifter_i3_LC_1_3_3 (
            .in0(N__5075),
            .in1(N__2075),
            .in2(N__2064),
            .in3(N__4915),
            .lcout(ctrl_idcodeArea_shifter_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4703),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_idcodeArea_shifter_i29_LC_1_3_4.C_ON=1'b0;
    defparam ctrl_idcodeArea_shifter_i29_LC_1_3_4.SEQ_MODE=4'b1000;
    defparam ctrl_idcodeArea_shifter_i29_LC_1_3_4.LUT_INIT=16'b1100000010001000;
    LogicCell40 ctrl_idcodeArea_shifter_i29_LC_1_3_4 (
            .in0(N__2049),
            .in1(N__4858),
            .in2(N__2349),
            .in3(N__5047),
            .lcout(ctrl_idcodeArea_shifter_29),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4703),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_idcodeArea_shifter_i30_LC_1_3_5.C_ON=1'b0;
    defparam ctrl_idcodeArea_shifter_i30_LC_1_3_5.SEQ_MODE=4'b1000;
    defparam ctrl_idcodeArea_shifter_i30_LC_1_3_5.LUT_INIT=16'b1101000010000000;
    LogicCell40 ctrl_idcodeArea_shifter_i30_LC_1_3_5 (
            .in0(N__5074),
            .in1(N__2048),
            .in2(N__4916),
            .in3(N__3717),
            .lcout(ctrl_idcodeArea_shifter_30),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4703),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_210_i4_4_lut_4_lut_LC_1_3_6.C_ON=1'b0;
    defparam mux_210_i4_4_lut_4_lut_LC_1_3_6.SEQ_MODE=4'b0000;
    defparam mux_210_i4_4_lut_4_lut_LC_1_3_6.LUT_INIT=16'b1110101001001010;
    LogicCell40 mux_210_i4_4_lut_4_lut_LC_1_3_6 (
            .in0(N__4053),
            .in1(N__4178),
            .in2(N__3973),
            .in3(N__3864),
            .lcout(n962),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_tap_fsm_state_3__I_0_i6_2_lut_LC_1_3_7.C_ON=1'b0;
    defparam ctrl_tap_fsm_state_3__I_0_i6_2_lut_LC_1_3_7.SEQ_MODE=4'b0000;
    defparam ctrl_tap_fsm_state_3__I_0_i6_2_lut_LC_1_3_7.LUT_INIT=16'b1100110011111111;
    LogicCell40 ctrl_tap_fsm_state_3__I_0_i6_2_lut_LC_1_3_7 (
            .in0(_gnd_net_),
            .in1(N__3658),
            .in2(_gnd_net_),
            .in3(N__4051),
            .lcout(n6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1073_2_lut_LC_1_4_0.C_ON=1'b0;
    defparam i1073_2_lut_LC_1_4_0.SEQ_MODE=4'b0000;
    defparam i1073_2_lut_LC_1_4_0.LUT_INIT=16'b1010101000000000;
    LogicCell40 i1073_2_lut_LC_1_4_0 (
            .in0(N__3962),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2106),
            .lcout(),
            .ltout(n1854_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1385_4_lut_LC_1_4_1.C_ON=1'b0;
    defparam i1385_4_lut_LC_1_4_1.SEQ_MODE=4'b0000;
    defparam i1385_4_lut_LC_1_4_1.LUT_INIT=16'b0000101011001100;
    LogicCell40 i1385_4_lut_LC_1_4_1 (
            .in0(N__2178),
            .in1(N__3780),
            .in2(N__2040),
            .in3(N__2751),
            .lcout(),
            .ltout(n2188_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_tap_fsm_state_i2_LC_1_4_2.C_ON=1'b0;
    defparam ctrl_tap_fsm_state_i2_LC_1_4_2.SEQ_MODE=4'b1000;
    defparam ctrl_tap_fsm_state_i2_LC_1_4_2.LUT_INIT=16'b0111010000110000;
    LogicCell40 ctrl_tap_fsm_state_i2_LC_1_4_2 (
            .in0(N__2753),
            .in1(N__2723),
            .in2(N__2133),
            .in3(N__2151),
            .lcout(ctrl_tap_fsm_state_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4701),
            .ce(),
            .sr(_gnd_net_));
    defparam i1431_2_lut_LC_1_4_3.C_ON=1'b0;
    defparam i1431_2_lut_LC_1_4_3.SEQ_MODE=4'b0000;
    defparam i1431_2_lut_LC_1_4_3.LUT_INIT=16'b1111111110101010;
    LogicCell40 i1431_2_lut_LC_1_4_3 (
            .in0(N__4182),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2750),
            .lcout(),
            .ltout(n2235_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_tap_fsm_state_i0_LC_1_4_4.C_ON=1'b0;
    defparam ctrl_tap_fsm_state_i0_LC_1_4_4.SEQ_MODE=4'b1000;
    defparam ctrl_tap_fsm_state_i0_LC_1_4_4.LUT_INIT=16'b0111111101001100;
    LogicCell40 ctrl_tap_fsm_state_i0_LC_1_4_4 (
            .in0(N__3961),
            .in1(N__2721),
            .in2(N__2130),
            .in3(N__2094),
            .lcout(ctrl_tap_fsm_state_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4701),
            .ce(),
            .sr(_gnd_net_));
    defparam i1427_2_lut_4_lut_LC_1_4_5.C_ON=1'b0;
    defparam i1427_2_lut_4_lut_LC_1_4_5.SEQ_MODE=4'b0000;
    defparam i1427_2_lut_4_lut_LC_1_4_5.LUT_INIT=16'b1100111011001100;
    LogicCell40 i1427_2_lut_4_lut_LC_1_4_5 (
            .in0(N__2160),
            .in1(N__3963),
            .in2(N__4213),
            .in3(N__3863),
            .lcout(),
            .ltout(n2202_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_tap_fsm_state_i1_LC_1_4_6.C_ON=1'b0;
    defparam ctrl_tap_fsm_state_i1_LC_1_4_6.SEQ_MODE=4'b1000;
    defparam ctrl_tap_fsm_state_i1_LC_1_4_6.LUT_INIT=16'b0111001101000000;
    LogicCell40 ctrl_tap_fsm_state_i1_LC_1_4_6 (
            .in0(N__2752),
            .in1(N__2722),
            .in2(N__2127),
            .in3(N__2463),
            .lcout(ctrl_tap_fsm_state_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4701),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_tap_fsm_state_i3_LC_1_4_7.C_ON=1'b0;
    defparam ctrl_tap_fsm_state_i3_LC_1_4_7.SEQ_MODE=4'b1000;
    defparam ctrl_tap_fsm_state_i3_LC_1_4_7.LUT_INIT=16'b0111001101100010;
    LogicCell40 ctrl_tap_fsm_state_i3_LC_1_4_7 (
            .in0(N__2724),
            .in1(N__2754),
            .in2(N__2124),
            .in3(N__2112),
            .lcout(ctrl_tap_fsm_state_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4701),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_3_lut_4_lut_LC_1_5_0.C_ON=1'b0;
    defparam i2_3_lut_4_lut_LC_1_5_0.SEQ_MODE=4'b0000;
    defparam i2_3_lut_4_lut_LC_1_5_0.LUT_INIT=16'b0000000000100000;
    LogicCell40 i2_3_lut_4_lut_LC_1_5_0 (
            .in0(N__4171),
            .in1(N__4063),
            .in2(N__3691),
            .in3(N__3854),
            .lcout(n1025),
            .ltout(n1025_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_209_i1_4_lut_LC_1_5_1.C_ON=1'b0;
    defparam mux_209_i1_4_lut_LC_1_5_1.SEQ_MODE=4'b0000;
    defparam mux_209_i1_4_lut_LC_1_5_1.LUT_INIT=16'b0000101001110111;
    LogicCell40 mux_209_i1_4_lut_LC_1_5_1 (
            .in0(N__3968),
            .in1(N__2184),
            .in2(N__2100),
            .in3(N__2177),
            .lcout(),
            .ltout(n960_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1391_3_lut_LC_1_5_2.C_ON=1'b0;
    defparam i1391_3_lut_LC_1_5_2.SEQ_MODE=4'b0000;
    defparam i1391_3_lut_LC_1_5_2.LUT_INIT=16'b1111000011001100;
    LogicCell40 i1391_3_lut_LC_1_5_2 (
            .in0(_gnd_net_),
            .in1(N__2166),
            .in2(N__2097),
            .in3(N__2748),
            .lcout(n2194),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i3_2_lut_3_lut_4_lut_LC_1_5_3.C_ON=1'b0;
    defparam i3_2_lut_3_lut_4_lut_LC_1_5_3.SEQ_MODE=4'b0000;
    defparam i3_2_lut_3_lut_4_lut_LC_1_5_3.LUT_INIT=16'b0000000000000010;
    LogicCell40 i3_2_lut_3_lut_4_lut_LC_1_5_3 (
            .in0(N__3855),
            .in1(N__4168),
            .in2(N__4083),
            .in3(N__3663),
            .lcout(n1023),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_4_lut_adj_2_LC_1_5_4.C_ON=1'b0;
    defparam i1_4_lut_4_lut_adj_2_LC_1_5_4.SEQ_MODE=4'b0000;
    defparam i1_4_lut_4_lut_adj_2_LC_1_5_4.LUT_INIT=16'b0000001000110000;
    LogicCell40 i1_4_lut_4_lut_adj_2_LC_1_5_4 (
            .in0(N__4169),
            .in1(N__4062),
            .in2(N__3690),
            .in3(N__3853),
            .lcout(n1027),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_210_i1_4_lut_LC_1_5_5.C_ON=1'b0;
    defparam mux_210_i1_4_lut_LC_1_5_5.SEQ_MODE=4'b0000;
    defparam mux_210_i1_4_lut_LC_1_5_5.LUT_INIT=16'b0000101000110000;
    LogicCell40 mux_210_i1_4_lut_LC_1_5_5 (
            .in0(N__3856),
            .in1(N__4170),
            .in2(N__3975),
            .in3(N__4068),
            .lcout(n965),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_LC_1_5_6.C_ON=1'b0;
    defparam i1_2_lut_LC_1_5_6.SEQ_MODE=4'b0000;
    defparam i1_2_lut_LC_1_5_6.LUT_INIT=16'b1010101000000000;
    LogicCell40 i1_2_lut_LC_1_5_6 (
            .in0(N__3670),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4064),
            .lcout(n5),
            .ltout(n5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1411_2_lut_4_lut_LC_1_5_7.C_ON=1'b0;
    defparam i1411_2_lut_4_lut_LC_1_5_7.SEQ_MODE=4'b0000;
    defparam i1411_2_lut_4_lut_LC_1_5_7.LUT_INIT=16'b1111111111011111;
    LogicCell40 i1411_2_lut_4_lut_LC_1_5_7 (
            .in0(N__3857),
            .in1(N__3972),
            .in2(N__2154),
            .in3(N__4172),
            .lcout(n2201),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam myClockArea_timeout_counter_value_313__i0_LC_1_6_0.C_ON=1'b1;
    defparam myClockArea_timeout_counter_value_313__i0_LC_1_6_0.SEQ_MODE=4'b1010;
    defparam myClockArea_timeout_counter_value_313__i0_LC_1_6_0.LUT_INIT=16'b1000001000101000;
    LogicCell40 myClockArea_timeout_counter_value_313__i0_LC_1_6_0 (
            .in0(N__2907),
            .in1(N__2664),
            .in2(_gnd_net_),
            .in3(N__2145),
            .lcout(myClockArea_timeout_counter_value_0),
            .ltout(),
            .carryin(bfn_1_6_0_),
            .carryout(n2009),
            .clk(N__5216),
            .ce(),
            .sr(N__3486));
    defparam myClockArea_timeout_counter_value_313__i1_LC_1_6_1.C_ON=1'b1;
    defparam myClockArea_timeout_counter_value_313__i1_LC_1_6_1.SEQ_MODE=4'b1010;
    defparam myClockArea_timeout_counter_value_313__i1_LC_1_6_1.LUT_INIT=16'b1000001000101000;
    LogicCell40 myClockArea_timeout_counter_value_313__i1_LC_1_6_1 (
            .in0(N__2877),
            .in1(N__2691),
            .in2(_gnd_net_),
            .in3(N__2142),
            .lcout(myClockArea_timeout_counter_value_1),
            .ltout(),
            .carryin(n2009),
            .carryout(n2010),
            .clk(N__5216),
            .ce(),
            .sr(N__3486));
    defparam myClockArea_timeout_counter_value_313__i2_LC_1_6_2.C_ON=1'b1;
    defparam myClockArea_timeout_counter_value_313__i2_LC_1_6_2.SEQ_MODE=4'b1010;
    defparam myClockArea_timeout_counter_value_313__i2_LC_1_6_2.LUT_INIT=16'b1000001000101000;
    LogicCell40 myClockArea_timeout_counter_value_313__i2_LC_1_6_2 (
            .in0(N__2908),
            .in1(N__2967),
            .in2(_gnd_net_),
            .in3(N__2139),
            .lcout(myClockArea_timeout_counter_value_2),
            .ltout(),
            .carryin(n2010),
            .carryout(n2011),
            .clk(N__5216),
            .ce(),
            .sr(N__3486));
    defparam myClockArea_timeout_counter_value_313__i3_LC_1_6_3.C_ON=1'b1;
    defparam myClockArea_timeout_counter_value_313__i3_LC_1_6_3.SEQ_MODE=4'b1010;
    defparam myClockArea_timeout_counter_value_313__i3_LC_1_6_3.LUT_INIT=16'b1000001000101000;
    LogicCell40 myClockArea_timeout_counter_value_313__i3_LC_1_6_3 (
            .in0(N__2878),
            .in1(N__2703),
            .in2(_gnd_net_),
            .in3(N__2136),
            .lcout(myClockArea_timeout_counter_value_3),
            .ltout(),
            .carryin(n2011),
            .carryout(n2012),
            .clk(N__5216),
            .ce(),
            .sr(N__3486));
    defparam myClockArea_timeout_counter_value_313__i4_LC_1_6_4.C_ON=1'b1;
    defparam myClockArea_timeout_counter_value_313__i4_LC_1_6_4.SEQ_MODE=4'b1010;
    defparam myClockArea_timeout_counter_value_313__i4_LC_1_6_4.LUT_INIT=16'b1000001000101000;
    LogicCell40 myClockArea_timeout_counter_value_313__i4_LC_1_6_4 (
            .in0(N__2909),
            .in1(N__3057),
            .in2(_gnd_net_),
            .in3(N__2211),
            .lcout(myClockArea_timeout_counter_value_4),
            .ltout(),
            .carryin(n2012),
            .carryout(n2013),
            .clk(N__5216),
            .ce(),
            .sr(N__3486));
    defparam myClockArea_timeout_counter_value_313__i5_LC_1_6_5.C_ON=1'b1;
    defparam myClockArea_timeout_counter_value_313__i5_LC_1_6_5.SEQ_MODE=4'b1010;
    defparam myClockArea_timeout_counter_value_313__i5_LC_1_6_5.LUT_INIT=16'b1000001000101000;
    LogicCell40 myClockArea_timeout_counter_value_313__i5_LC_1_6_5 (
            .in0(N__2879),
            .in1(N__2678),
            .in2(_gnd_net_),
            .in3(N__2208),
            .lcout(myClockArea_timeout_counter_value_5),
            .ltout(),
            .carryin(n2013),
            .carryout(n2014),
            .clk(N__5216),
            .ce(),
            .sr(N__3486));
    defparam myClockArea_timeout_counter_value_313__i6_LC_1_6_6.C_ON=1'b1;
    defparam myClockArea_timeout_counter_value_313__i6_LC_1_6_6.SEQ_MODE=4'b1010;
    defparam myClockArea_timeout_counter_value_313__i6_LC_1_6_6.LUT_INIT=16'b1000001000101000;
    LogicCell40 myClockArea_timeout_counter_value_313__i6_LC_1_6_6 (
            .in0(N__2910),
            .in1(N__3045),
            .in2(_gnd_net_),
            .in3(N__2205),
            .lcout(myClockArea_timeout_counter_value_6),
            .ltout(),
            .carryin(n2014),
            .carryout(n2015),
            .clk(N__5216),
            .ce(),
            .sr(N__3486));
    defparam myClockArea_timeout_counter_value_313__i7_LC_1_6_7.C_ON=1'b1;
    defparam myClockArea_timeout_counter_value_313__i7_LC_1_6_7.SEQ_MODE=4'b1010;
    defparam myClockArea_timeout_counter_value_313__i7_LC_1_6_7.LUT_INIT=16'b1000001000101000;
    LogicCell40 myClockArea_timeout_counter_value_313__i7_LC_1_6_7 (
            .in0(N__2880),
            .in1(N__2583),
            .in2(_gnd_net_),
            .in3(N__2202),
            .lcout(myClockArea_timeout_counter_value_7),
            .ltout(),
            .carryin(n2015),
            .carryout(n2016),
            .clk(N__5216),
            .ce(),
            .sr(N__3486));
    defparam myClockArea_timeout_counter_value_313__i8_LC_1_7_0.C_ON=1'b1;
    defparam myClockArea_timeout_counter_value_313__i8_LC_1_7_0.SEQ_MODE=4'b1010;
    defparam myClockArea_timeout_counter_value_313__i8_LC_1_7_0.LUT_INIT=16'b1000001000101000;
    LogicCell40 myClockArea_timeout_counter_value_313__i8_LC_1_7_0 (
            .in0(N__2906),
            .in1(N__2994),
            .in2(_gnd_net_),
            .in3(N__2199),
            .lcout(myClockArea_timeout_counter_value_8),
            .ltout(),
            .carryin(bfn_1_7_0_),
            .carryout(n2017),
            .clk(N__5215),
            .ce(),
            .sr(N__3463));
    defparam myClockArea_timeout_counter_value_313__i9_LC_1_7_1.C_ON=1'b1;
    defparam myClockArea_timeout_counter_value_313__i9_LC_1_7_1.SEQ_MODE=4'b1010;
    defparam myClockArea_timeout_counter_value_313__i9_LC_1_7_1.LUT_INIT=16'b1000001000101000;
    LogicCell40 myClockArea_timeout_counter_value_313__i9_LC_1_7_1 (
            .in0(N__2873),
            .in1(N__2652),
            .in2(_gnd_net_),
            .in3(N__2196),
            .lcout(myClockArea_timeout_counter_value_9),
            .ltout(),
            .carryin(n2017),
            .carryout(n2018),
            .clk(N__5215),
            .ce(),
            .sr(N__3463));
    defparam myClockArea_timeout_counter_value_313__i10_LC_1_7_2.C_ON=1'b1;
    defparam myClockArea_timeout_counter_value_313__i10_LC_1_7_2.SEQ_MODE=4'b1010;
    defparam myClockArea_timeout_counter_value_313__i10_LC_1_7_2.LUT_INIT=16'b1000001000101000;
    LogicCell40 myClockArea_timeout_counter_value_313__i10_LC_1_7_2 (
            .in0(N__2903),
            .in1(N__2981),
            .in2(_gnd_net_),
            .in3(N__2193),
            .lcout(myClockArea_timeout_counter_value_10),
            .ltout(),
            .carryin(n2018),
            .carryout(n2019),
            .clk(N__5215),
            .ce(),
            .sr(N__3463));
    defparam myClockArea_timeout_counter_value_313__i11_LC_1_7_3.C_ON=1'b1;
    defparam myClockArea_timeout_counter_value_313__i11_LC_1_7_3.SEQ_MODE=4'b1010;
    defparam myClockArea_timeout_counter_value_313__i11_LC_1_7_3.LUT_INIT=16'b1000001000101000;
    LogicCell40 myClockArea_timeout_counter_value_313__i11_LC_1_7_3 (
            .in0(N__2870),
            .in1(N__2778),
            .in2(_gnd_net_),
            .in3(N__2190),
            .lcout(myClockArea_timeout_counter_value_11),
            .ltout(),
            .carryin(n2019),
            .carryout(n2020),
            .clk(N__5215),
            .ce(),
            .sr(N__3463));
    defparam myClockArea_timeout_counter_value_313__i12_LC_1_7_4.C_ON=1'b1;
    defparam myClockArea_timeout_counter_value_313__i12_LC_1_7_4.SEQ_MODE=4'b1010;
    defparam myClockArea_timeout_counter_value_313__i12_LC_1_7_4.LUT_INIT=16'b1000001000101000;
    LogicCell40 myClockArea_timeout_counter_value_313__i12_LC_1_7_4 (
            .in0(N__2904),
            .in1(N__2624),
            .in2(_gnd_net_),
            .in3(N__2187),
            .lcout(myClockArea_timeout_counter_value_12),
            .ltout(),
            .carryin(n2020),
            .carryout(n2021),
            .clk(N__5215),
            .ce(),
            .sr(N__3463));
    defparam myClockArea_timeout_counter_value_313__i13_LC_1_7_5.C_ON=1'b1;
    defparam myClockArea_timeout_counter_value_313__i13_LC_1_7_5.SEQ_MODE=4'b1010;
    defparam myClockArea_timeout_counter_value_313__i13_LC_1_7_5.LUT_INIT=16'b1000001000101000;
    LogicCell40 myClockArea_timeout_counter_value_313__i13_LC_1_7_5 (
            .in0(N__2871),
            .in1(N__2940),
            .in2(_gnd_net_),
            .in3(N__2238),
            .lcout(myClockArea_timeout_counter_value_13),
            .ltout(),
            .carryin(n2021),
            .carryout(n2022),
            .clk(N__5215),
            .ce(),
            .sr(N__3463));
    defparam myClockArea_timeout_counter_value_313__i14_LC_1_7_6.C_ON=1'b1;
    defparam myClockArea_timeout_counter_value_313__i14_LC_1_7_6.SEQ_MODE=4'b1010;
    defparam myClockArea_timeout_counter_value_313__i14_LC_1_7_6.LUT_INIT=16'b1000001000101000;
    LogicCell40 myClockArea_timeout_counter_value_313__i14_LC_1_7_6 (
            .in0(N__2905),
            .in1(N__2610),
            .in2(_gnd_net_),
            .in3(N__2235),
            .lcout(myClockArea_timeout_counter_value_14),
            .ltout(),
            .carryin(n2022),
            .carryout(n2023),
            .clk(N__5215),
            .ce(),
            .sr(N__3463));
    defparam myClockArea_timeout_counter_value_313__i15_LC_1_7_7.C_ON=1'b1;
    defparam myClockArea_timeout_counter_value_313__i15_LC_1_7_7.SEQ_MODE=4'b1010;
    defparam myClockArea_timeout_counter_value_313__i15_LC_1_7_7.LUT_INIT=16'b1000001000101000;
    LogicCell40 myClockArea_timeout_counter_value_313__i15_LC_1_7_7 (
            .in0(N__2872),
            .in1(N__2805),
            .in2(_gnd_net_),
            .in3(N__2232),
            .lcout(myClockArea_timeout_counter_value_15),
            .ltout(),
            .carryin(n2023),
            .carryout(n2024),
            .clk(N__5215),
            .ce(),
            .sr(N__3463));
    defparam myClockArea_timeout_counter_value_313__i16_LC_1_8_0.C_ON=1'b1;
    defparam myClockArea_timeout_counter_value_313__i16_LC_1_8_0.SEQ_MODE=4'b1010;
    defparam myClockArea_timeout_counter_value_313__i16_LC_1_8_0.LUT_INIT=16'b1000001000101000;
    LogicCell40 myClockArea_timeout_counter_value_313__i16_LC_1_8_0 (
            .in0(N__2899),
            .in1(N__3018),
            .in2(_gnd_net_),
            .in3(N__2229),
            .lcout(myClockArea_timeout_counter_value_16),
            .ltout(),
            .carryin(bfn_1_8_0_),
            .carryout(n2025),
            .clk(N__5213),
            .ce(),
            .sr(N__3478));
    defparam myClockArea_timeout_counter_value_313__i17_LC_1_8_1.C_ON=1'b1;
    defparam myClockArea_timeout_counter_value_313__i17_LC_1_8_1.SEQ_MODE=4'b1010;
    defparam myClockArea_timeout_counter_value_313__i17_LC_1_8_1.LUT_INIT=16'b1000001000101000;
    LogicCell40 myClockArea_timeout_counter_value_313__i17_LC_1_8_1 (
            .in0(N__2874),
            .in1(N__3006),
            .in2(_gnd_net_),
            .in3(N__2226),
            .lcout(myClockArea_timeout_counter_value_17),
            .ltout(),
            .carryin(n2025),
            .carryout(n2026),
            .clk(N__5213),
            .ce(),
            .sr(N__3478));
    defparam myClockArea_timeout_counter_value_313__i18_LC_1_8_2.C_ON=1'b1;
    defparam myClockArea_timeout_counter_value_313__i18_LC_1_8_2.SEQ_MODE=4'b1010;
    defparam myClockArea_timeout_counter_value_313__i18_LC_1_8_2.LUT_INIT=16'b1000001000101000;
    LogicCell40 myClockArea_timeout_counter_value_313__i18_LC_1_8_2 (
            .in0(N__2900),
            .in1(N__2639),
            .in2(_gnd_net_),
            .in3(N__2223),
            .lcout(myClockArea_timeout_counter_value_18),
            .ltout(),
            .carryin(n2026),
            .carryout(n2027),
            .clk(N__5213),
            .ce(),
            .sr(N__3478));
    defparam myClockArea_timeout_counter_value_313__i19_LC_1_8_3.C_ON=1'b1;
    defparam myClockArea_timeout_counter_value_313__i19_LC_1_8_3.SEQ_MODE=4'b1010;
    defparam myClockArea_timeout_counter_value_313__i19_LC_1_8_3.LUT_INIT=16'b1000001000101000;
    LogicCell40 myClockArea_timeout_counter_value_313__i19_LC_1_8_3 (
            .in0(N__2875),
            .in1(N__2817),
            .in2(_gnd_net_),
            .in3(N__2220),
            .lcout(myClockArea_timeout_counter_value_19),
            .ltout(),
            .carryin(n2027),
            .carryout(n2028),
            .clk(N__5213),
            .ce(),
            .sr(N__3478));
    defparam myClockArea_timeout_counter_value_313__i20_LC_1_8_4.C_ON=1'b1;
    defparam myClockArea_timeout_counter_value_313__i20_LC_1_8_4.SEQ_MODE=4'b1010;
    defparam myClockArea_timeout_counter_value_313__i20_LC_1_8_4.LUT_INIT=16'b1000001000101000;
    LogicCell40 myClockArea_timeout_counter_value_313__i20_LC_1_8_4 (
            .in0(N__2901),
            .in1(N__2792),
            .in2(_gnd_net_),
            .in3(N__2217),
            .lcout(myClockArea_timeout_counter_value_20),
            .ltout(),
            .carryin(n2028),
            .carryout(n2029),
            .clk(N__5213),
            .ce(),
            .sr(N__3478));
    defparam myClockArea_timeout_counter_value_313__i21_LC_1_8_5.C_ON=1'b1;
    defparam myClockArea_timeout_counter_value_313__i21_LC_1_8_5.SEQ_MODE=4'b1010;
    defparam myClockArea_timeout_counter_value_313__i21_LC_1_8_5.LUT_INIT=16'b1000001000101000;
    LogicCell40 myClockArea_timeout_counter_value_313__i21_LC_1_8_5 (
            .in0(N__2876),
            .in1(N__2570),
            .in2(_gnd_net_),
            .in3(N__2214),
            .lcout(myClockArea_timeout_counter_value_21),
            .ltout(),
            .carryin(n2029),
            .carryout(n2030),
            .clk(N__5213),
            .ce(),
            .sr(N__3478));
    defparam myClockArea_timeout_counter_value_313__i22_LC_1_8_6.C_ON=1'b0;
    defparam myClockArea_timeout_counter_value_313__i22_LC_1_8_6.SEQ_MODE=4'b1010;
    defparam myClockArea_timeout_counter_value_313__i22_LC_1_8_6.LUT_INIT=16'b1000001000101000;
    LogicCell40 myClockArea_timeout_counter_value_313__i22_LC_1_8_6 (
            .in0(N__2902),
            .in1(N__3032),
            .in2(_gnd_net_),
            .in3(N__2298),
            .lcout(myClockArea_timeout_counter_value_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5213),
            .ce(),
            .sr(N__3478));
    defparam ctrl_tap_instruction_i4_LC_2_1_0.C_ON=1'b0;
    defparam ctrl_tap_instruction_i4_LC_2_1_0.SEQ_MODE=4'b1000;
    defparam ctrl_tap_instruction_i4_LC_2_1_0.LUT_INIT=16'b1100100001000000;
    LogicCell40 ctrl_tap_instruction_i4_LC_2_1_0 (
            .in0(N__2265),
            .in1(N__4927),
            .in2(N__3273),
            .in3(N__3360),
            .lcout(ctrl_tap_instruction_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4710),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_tap_instruction_i0_LC_2_1_1.C_ON=1'b0;
    defparam ctrl_tap_instruction_i0_LC_2_1_1.SEQ_MODE=4'b1000;
    defparam ctrl_tap_instruction_i0_LC_2_1_1.LUT_INIT=16'b1000100010100000;
    LogicCell40 ctrl_tap_instruction_i0_LC_2_1_1 (
            .in0(N__4923),
            .in1(N__3128),
            .in2(N__3099),
            .in3(N__2268),
            .lcout(ctrl_tap_instruction_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4710),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_8_LC_2_1_2.C_ON=1'b0;
    defparam i1_2_lut_adj_8_LC_2_1_2.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_8_LC_2_1_2.LUT_INIT=16'b1111111111001100;
    LogicCell40 i1_2_lut_adj_8_LC_2_1_2 (
            .in0(_gnd_net_),
            .in1(N__4341),
            .in2(_gnd_net_),
            .in3(N__2295),
            .lcout(),
            .ltout(n4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i395_4_lut_LC_2_1_3.C_ON=1'b0;
    defparam i395_4_lut_LC_2_1_3.SEQ_MODE=4'b0000;
    defparam i395_4_lut_LC_2_1_3.LUT_INIT=16'b1111111000000010;
    LogicCell40 i395_4_lut_LC_2_1_3 (
            .in0(N__2364),
            .in1(N__2423),
            .in2(N__2289),
            .in3(N__2388),
            .lcout(),
            .ltout(ctrl_tap_tdoUnbufferd_N_223_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i398_4_lut_LC_2_1_4.C_ON=1'b0;
    defparam i398_4_lut_LC_2_1_4.SEQ_MODE=4'b0000;
    defparam i398_4_lut_LC_2_1_4.LUT_INIT=16'b1111000011100010;
    LogicCell40 i398_4_lut_LC_2_1_4 (
            .in0(N__3509),
            .in1(N__3761),
            .in2(N__2286),
            .in3(N__4342),
            .lcout(ctrl_tap_tdoUnbufferd),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_tap_instruction_i3_LC_2_1_5.C_ON=1'b0;
    defparam ctrl_tap_instruction_i3_LC_2_1_5.SEQ_MODE=4'b1000;
    defparam ctrl_tap_instruction_i3_LC_2_1_5.LUT_INIT=16'b1010100000100000;
    LogicCell40 ctrl_tap_instruction_i3_LC_2_1_5 (
            .in0(N__4924),
            .in1(N__2266),
            .in2(N__3225),
            .in3(N__3247),
            .lcout(ctrl_tap_instruction_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4710),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_tap_instruction_i2_LC_2_1_6.C_ON=1'b0;
    defparam ctrl_tap_instruction_i2_LC_2_1_6.SEQ_MODE=4'b1000;
    defparam ctrl_tap_instruction_i2_LC_2_1_6.LUT_INIT=16'b1111011110110011;
    LogicCell40 ctrl_tap_instruction_i2_LC_2_1_6 (
            .in0(N__2264),
            .in1(N__4926),
            .in2(N__3405),
            .in3(N__3375),
            .lcout(ctrl_tap_instruction_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4710),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_tap_instruction_i7_LC_2_1_7.C_ON=1'b0;
    defparam ctrl_tap_instruction_i7_LC_2_1_7.SEQ_MODE=4'b1000;
    defparam ctrl_tap_instruction_i7_LC_2_1_7.LUT_INIT=16'b1010000010001000;
    LogicCell40 ctrl_tap_instruction_i7_LC_2_1_7 (
            .in0(N__4925),
            .in1(N__3207),
            .in2(N__3300),
            .in3(N__2267),
            .lcout(ctrl_tap_instruction_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4710),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_LC_2_2_0.C_ON=1'b0;
    defparam i1_2_lut_3_lut_LC_2_2_0.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_LC_2_2_0.LUT_INIT=16'b1111111111101110;
    LogicCell40 i1_2_lut_3_lut_LC_2_2_0 (
            .in0(N__4183),
            .in1(N__4072),
            .in2(_gnd_net_),
            .in3(N__3868),
            .lcout(),
            .ltout(n1313_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_tap_bypass_I_0_4_lut_LC_2_2_1.C_ON=1'b0;
    defparam ctrl_tap_bypass_I_0_4_lut_LC_2_2_1.SEQ_MODE=4'b0000;
    defparam ctrl_tap_bypass_I_0_4_lut_LC_2_2_1.LUT_INIT=16'b1010110010101010;
    LogicCell40 ctrl_tap_bypass_I_0_4_lut_LC_2_2_1 (
            .in0(N__5157),
            .in1(N__3092),
            .in2(N__2391),
            .in3(N__3682),
            .lcout(ctrl_tap_tdoUnbufferd_N_224),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_idcodeArea_shifter_i25_LC_2_2_2.C_ON=1'b0;
    defparam ctrl_idcodeArea_shifter_i25_LC_2_2_2.SEQ_MODE=4'b1000;
    defparam ctrl_idcodeArea_shifter_i25_LC_2_2_2.LUT_INIT=16'b1101100011111111;
    LogicCell40 ctrl_idcodeArea_shifter_i25_LC_2_2_2 (
            .in0(N__5039),
            .in1(N__2456),
            .in2(N__2310),
            .in3(N__4857),
            .lcout(ctrl_idcodeArea_shifter_25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4708),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_idcodeArea_shifter_i0_LC_2_2_3.C_ON=1'b0;
    defparam ctrl_idcodeArea_shifter_i0_LC_2_2_3.SEQ_MODE=4'b1000;
    defparam ctrl_idcodeArea_shifter_i0_LC_2_2_3.LUT_INIT=16'b1111110101110101;
    LogicCell40 ctrl_idcodeArea_shifter_i0_LC_2_2_3 (
            .in0(N__4854),
            .in1(N__5041),
            .in2(N__2382),
            .in3(N__2363),
            .lcout(ctrl_idcodeArea_shifter_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4708),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_9_LC_2_2_4.C_ON=1'b0;
    defparam i1_2_lut_adj_9_LC_2_2_4.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_9_LC_2_2_4.LUT_INIT=16'b1111111111001100;
    LogicCell40 i1_2_lut_adj_9_LC_2_2_4 (
            .in0(_gnd_net_),
            .in1(N__3125),
            .in2(_gnd_net_),
            .in3(N__3428),
            .lcout(n2119),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_idcodeArea_shifter_i28_LC_2_2_5.C_ON=1'b0;
    defparam ctrl_idcodeArea_shifter_i28_LC_2_2_5.SEQ_MODE=4'b1000;
    defparam ctrl_idcodeArea_shifter_i28_LC_2_2_5.LUT_INIT=16'b1010000010001000;
    LogicCell40 ctrl_idcodeArea_shifter_i28_LC_2_2_5 (
            .in0(N__4856),
            .in1(N__2348),
            .in2(N__2334),
            .in3(N__5043),
            .lcout(ctrl_idcodeArea_shifter_28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4708),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_idcodeArea_shifter_i27_LC_2_2_6.C_ON=1'b0;
    defparam ctrl_idcodeArea_shifter_i27_LC_2_2_6.SEQ_MODE=4'b1000;
    defparam ctrl_idcodeArea_shifter_i27_LC_2_2_6.LUT_INIT=16'b1101000010000000;
    LogicCell40 ctrl_idcodeArea_shifter_i27_LC_2_2_6 (
            .in0(N__5040),
            .in1(N__2318),
            .in2(N__4919),
            .in3(N__2330),
            .lcout(ctrl_idcodeArea_shifter_27),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4708),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_idcodeArea_shifter_i26_LC_2_2_7.C_ON=1'b0;
    defparam ctrl_idcodeArea_shifter_i26_LC_2_2_7.SEQ_MODE=4'b1000;
    defparam ctrl_idcodeArea_shifter_i26_LC_2_2_7.LUT_INIT=16'b1101110111110101;
    LogicCell40 ctrl_idcodeArea_shifter_i26_LC_2_2_7 (
            .in0(N__4855),
            .in1(N__2306),
            .in2(N__2322),
            .in3(N__5042),
            .lcout(ctrl_idcodeArea_shifter_26),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4708),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_idcodeArea_shifter_i22_LC_2_3_0.C_ON=1'b0;
    defparam ctrl_idcodeArea_shifter_i22_LC_2_3_0.SEQ_MODE=4'b1000;
    defparam ctrl_idcodeArea_shifter_i22_LC_2_3_0.LUT_INIT=16'b1010111111001111;
    LogicCell40 ctrl_idcodeArea_shifter_i22_LC_2_3_0 (
            .in0(N__3566),
            .in1(N__2400),
            .in2(N__4918),
            .in3(N__5038),
            .lcout(ctrl_idcodeArea_shifter_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4706),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_tap_fsm_state_3__I_0_i7_2_lut_4_lut_LC_2_3_1.C_ON=1'b0;
    defparam ctrl_tap_fsm_state_3__I_0_i7_2_lut_4_lut_LC_2_3_1.SEQ_MODE=4'b0000;
    defparam ctrl_tap_fsm_state_3__I_0_i7_2_lut_4_lut_LC_2_3_1.LUT_INIT=16'b1111011111111111;
    LogicCell40 ctrl_tap_fsm_state_3__I_0_i7_2_lut_4_lut_LC_2_3_1 (
            .in0(N__4146),
            .in1(N__4038),
            .in2(N__3681),
            .in3(N__3838),
            .lcout(n7_adj_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_ledsArea_store_i0_i5_LC_2_3_2.C_ON=1'b0;
    defparam ctrl_ledsArea_store_i0_i5_LC_2_3_2.SEQ_MODE=4'b1000;
    defparam ctrl_ledsArea_store_i0_i5_LC_2_3_2.LUT_INIT=16'b1110111001000100;
    LogicCell40 ctrl_ledsArea_store_i0_i5_LC_2_3_2 (
            .in0(N__2509),
            .in1(N__4485),
            .in2(_gnd_net_),
            .in3(N__4496),
            .lcout(ctrl_ledsArea_store_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4706),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_idcodeArea_shifter_i24_LC_2_3_3.C_ON=1'b0;
    defparam ctrl_idcodeArea_shifter_i24_LC_2_3_3.SEQ_MODE=4'b1000;
    defparam ctrl_idcodeArea_shifter_i24_LC_2_3_3.LUT_INIT=16'b1110111101001111;
    LogicCell40 ctrl_idcodeArea_shifter_i24_LC_2_3_3 (
            .in0(N__5037),
            .in1(N__2457),
            .in2(N__4917),
            .in3(N__2412),
            .lcout(ctrl_idcodeArea_shifter_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4706),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_4_lut_adj_7_LC_2_3_4.C_ON=1'b0;
    defparam i1_2_lut_3_lut_4_lut_adj_7_LC_2_3_4.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_4_lut_adj_7_LC_2_3_4.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_2_lut_3_lut_4_lut_adj_7_LC_2_3_4 (
            .in0(N__3839),
            .in1(N__4147),
            .in2(N__4071),
            .in3(N__3649),
            .lcout(n1582),
            .ltout(n1582_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1375_4_lut_LC_2_3_5.C_ON=1'b0;
    defparam i1375_4_lut_LC_2_3_5.SEQ_MODE=4'b0000;
    defparam i1375_4_lut_LC_2_3_5.LUT_INIT=16'b1111000011100000;
    LogicCell40 i1375_4_lut_LC_2_3_5 (
            .in0(N__2445),
            .in1(N__2439),
            .in2(N__2427),
            .in3(N__2424),
            .lcout(n2178),
            .ltout(n2178_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_idcodeArea_shifter_i23_LC_2_3_6.C_ON=1'b0;
    defparam ctrl_idcodeArea_shifter_i23_LC_2_3_6.SEQ_MODE=4'b1000;
    defparam ctrl_idcodeArea_shifter_i23_LC_2_3_6.LUT_INIT=16'b1100101000000000;
    LogicCell40 ctrl_idcodeArea_shifter_i23_LC_2_3_6 (
            .in0(N__2411),
            .in1(N__2399),
            .in2(N__2403),
            .in3(N__4870),
            .lcout(ctrl_idcodeArea_shifter_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4706),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_ledsArea_store_i0_i1_LC_2_3_7.C_ON=1'b0;
    defparam ctrl_ledsArea_store_i0_i1_LC_2_3_7.SEQ_MODE=4'b1000;
    defparam ctrl_ledsArea_store_i0_i1_LC_2_3_7.LUT_INIT=16'b1011101110001000;
    LogicCell40 ctrl_ledsArea_store_i0_i1_LC_2_3_7 (
            .in0(N__3532),
            .in1(N__2508),
            .in2(_gnd_net_),
            .in3(N__3510),
            .lcout(io_leds_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4706),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_idcodeArea_shifter_i7_LC_2_4_0.C_ON=1'b0;
    defparam ctrl_idcodeArea_shifter_i7_LC_2_4_0.SEQ_MODE=4'b1000;
    defparam ctrl_idcodeArea_shifter_i7_LC_2_4_0.LUT_INIT=16'b1100000010001000;
    LogicCell40 ctrl_idcodeArea_shifter_i7_LC_2_4_0 (
            .in0(N__2486),
            .in1(N__4864),
            .in2(N__2541),
            .in3(N__5046),
            .lcout(ctrl_idcodeArea_shifter_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4704),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_ledsArea_store_i0_i3_LC_2_4_1.C_ON=1'b0;
    defparam ctrl_ledsArea_store_i0_i3_LC_2_4_1.SEQ_MODE=4'b1000;
    defparam ctrl_ledsArea_store_i0_i3_LC_2_4_1.LUT_INIT=16'b1110111001000100;
    LogicCell40 ctrl_ledsArea_store_i0_i3_LC_2_4_1 (
            .in0(N__2511),
            .in1(N__4575),
            .in2(_gnd_net_),
            .in3(N__4588),
            .lcout(io_leds_c_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4704),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_ledsArea_store_i0_i2_LC_2_4_2.C_ON=1'b0;
    defparam ctrl_ledsArea_store_i0_i2_LC_2_4_2.SEQ_MODE=4'b1000;
    defparam ctrl_ledsArea_store_i0_i2_LC_2_4_2.LUT_INIT=16'b1100110010101010;
    LogicCell40 ctrl_ledsArea_store_i0_i2_LC_2_4_2 (
            .in0(N__4623),
            .in1(N__4636),
            .in2(_gnd_net_),
            .in3(N__2510),
            .lcout(io_leds_c_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4704),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_ledsArea_store_i0_i4_LC_2_4_3.C_ON=1'b0;
    defparam ctrl_ledsArea_store_i0_i4_LC_2_4_3.SEQ_MODE=4'b1000;
    defparam ctrl_ledsArea_store_i0_i4_LC_2_4_3.LUT_INIT=16'b1111101001010000;
    LogicCell40 ctrl_ledsArea_store_i0_i4_LC_2_4_3 (
            .in0(N__2512),
            .in1(_gnd_net_),
            .in2(N__4524),
            .in3(N__4537),
            .lcout(io_leds_c_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4704),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_idcodeArea_shifter_i5_LC_2_4_4.C_ON=1'b0;
    defparam ctrl_idcodeArea_shifter_i5_LC_2_4_4.SEQ_MODE=4'b1000;
    defparam ctrl_idcodeArea_shifter_i5_LC_2_4_4.LUT_INIT=16'b1111001110111011;
    LogicCell40 ctrl_idcodeArea_shifter_i5_LC_2_4_4 (
            .in0(N__2528),
            .in1(N__4863),
            .in2(N__2556),
            .in3(N__5045),
            .lcout(ctrl_idcodeArea_shifter_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4704),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_idcodeArea_shifter_i6_LC_2_4_5.C_ON=1'b0;
    defparam ctrl_idcodeArea_shifter_i6_LC_2_4_5.SEQ_MODE=4'b1000;
    defparam ctrl_idcodeArea_shifter_i6_LC_2_4_5.LUT_INIT=16'b1110010000000000;
    LogicCell40 ctrl_idcodeArea_shifter_i6_LC_2_4_5 (
            .in0(N__5044),
            .in1(N__2540),
            .in2(N__2529),
            .in3(N__4877),
            .lcout(ctrl_idcodeArea_shifter_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4704),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_ledsArea_store_i0_i8_LC_2_4_6.C_ON=1'b0;
    defparam ctrl_ledsArea_store_i0_i8_LC_2_4_6.SEQ_MODE=4'b1000;
    defparam ctrl_ledsArea_store_i0_i8_LC_2_4_6.LUT_INIT=16'b1100110010101010;
    LogicCell40 ctrl_ledsArea_store_i0_i8_LC_2_4_6 (
            .in0(N__4254),
            .in1(N__4306),
            .in2(_gnd_net_),
            .in3(N__2514),
            .lcout(io_leds_c_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4704),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_ledsArea_store_i0_i6_LC_2_4_7.C_ON=1'b0;
    defparam ctrl_ledsArea_store_i0_i6_LC_2_4_7.SEQ_MODE=4'b1000;
    defparam ctrl_ledsArea_store_i0_i6_LC_2_4_7.LUT_INIT=16'b1111101001010000;
    LogicCell40 ctrl_ledsArea_store_i0_i6_LC_2_4_7 (
            .in0(N__2513),
            .in1(_gnd_net_),
            .in2(N__4434),
            .in3(N__4450),
            .lcout(io_leds_c_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4704),
            .ce(),
            .sr(_gnd_net_));
    defparam i1337_2_lut_LC_2_5_0.C_ON=1'b0;
    defparam i1337_2_lut_LC_2_5_0.SEQ_MODE=4'b0000;
    defparam i1337_2_lut_LC_2_5_0.LUT_INIT=16'b1111111111001100;
    LogicCell40 i1337_2_lut_LC_2_5_0 (
            .in0(_gnd_net_),
            .in1(N__3964),
            .in2(_gnd_net_),
            .in3(N__4065),
            .lcout(n2140),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_idcodeArea_shifter_i8_LC_2_5_1.C_ON=1'b0;
    defparam ctrl_idcodeArea_shifter_i8_LC_2_5_1.SEQ_MODE=4'b1000;
    defparam ctrl_idcodeArea_shifter_i8_LC_2_5_1.LUT_INIT=16'b1111001110111011;
    LogicCell40 ctrl_idcodeArea_shifter_i8_LC_2_5_1 (
            .in0(N__2597),
            .in1(N__4899),
            .in2(N__2487),
            .in3(N__5064),
            .lcout(ctrl_idcodeArea_shifter_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4702),
            .ce(),
            .sr(_gnd_net_));
    defparam i20_4_lut_3_lut_LC_2_5_2.C_ON=1'b0;
    defparam i20_4_lut_3_lut_LC_2_5_2.SEQ_MODE=4'b0000;
    defparam i20_4_lut_3_lut_LC_2_5_2.LUT_INIT=16'b0001000110001000;
    LogicCell40 i20_4_lut_3_lut_LC_2_5_2 (
            .in0(N__4176),
            .in1(N__3677),
            .in2(_gnd_net_),
            .in3(N__3858),
            .lcout(),
            .ltout(n9_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1388_4_lut_LC_2_5_3.C_ON=1'b0;
    defparam i1388_4_lut_LC_2_5_3.SEQ_MODE=4'b0000;
    defparam i1388_4_lut_LC_2_5_3.LUT_INIT=16'b0101000000110011;
    LogicCell40 i1388_4_lut_LC_2_5_3 (
            .in0(N__2472),
            .in1(N__2709),
            .in2(N__2466),
            .in3(N__2749),
            .lcout(n2191),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_LC_2_5_4.C_ON=1'b0;
    defparam i1_4_lut_LC_2_5_4.SEQ_MODE=4'b0000;
    defparam i1_4_lut_LC_2_5_4.LUT_INIT=16'b1000001100110111;
    LogicCell40 i1_4_lut_LC_2_5_4 (
            .in0(N__4173),
            .in1(N__4066),
            .in2(N__3692),
            .in3(N__3859),
            .lcout(n12_adj_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i988_4_lut_4_lut_LC_2_5_5.C_ON=1'b0;
    defparam i988_4_lut_4_lut_LC_2_5_5.SEQ_MODE=4'b0000;
    defparam i988_4_lut_4_lut_LC_2_5_5.LUT_INIT=16'b0111000000000001;
    LogicCell40 i988_4_lut_4_lut_LC_2_5_5 (
            .in0(N__3861),
            .in1(N__4177),
            .in2(N__3694),
            .in3(N__4070),
            .lcout(n1769),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_4_lut_LC_2_5_6.C_ON=1'b0;
    defparam i1_2_lut_3_lut_4_lut_LC_2_5_6.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_4_lut_LC_2_5_6.LUT_INIT=16'b1111101111111111;
    LogicCell40 i1_2_lut_3_lut_4_lut_LC_2_5_6 (
            .in0(N__4175),
            .in1(N__4067),
            .in2(N__3693),
            .in3(N__3862),
            .lcout(n7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_210_i2_4_lut_LC_2_5_7.C_ON=1'b0;
    defparam mux_210_i2_4_lut_LC_2_5_7.SEQ_MODE=4'b0000;
    defparam mux_210_i2_4_lut_LC_2_5_7.LUT_INIT=16'b1010000011001100;
    LogicCell40 mux_210_i2_4_lut_LC_2_5_7 (
            .in0(N__3860),
            .in1(N__4174),
            .in2(N__3974),
            .in3(N__4069),
            .lcout(n1864),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1361_4_lut_LC_2_6_0.C_ON=1'b0;
    defparam i1361_4_lut_LC_2_6_0.SEQ_MODE=4'b0000;
    defparam i1361_4_lut_LC_2_6_0.LUT_INIT=16'b1000000000000000;
    LogicCell40 i1361_4_lut_LC_2_6_0 (
            .in0(N__2702),
            .in1(N__2690),
            .in2(N__2679),
            .in3(N__2663),
            .lcout(n2164),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i5_4_lut_adj_3_LC_2_6_2.C_ON=1'b0;
    defparam i5_4_lut_adj_3_LC_2_6_2.SEQ_MODE=4'b0000;
    defparam i5_4_lut_adj_3_LC_2_6_2.LUT_INIT=16'b1111111111111110;
    LogicCell40 i5_4_lut_adj_3_LC_2_6_2 (
            .in0(N__2651),
            .in1(N__2640),
            .in2(N__2625),
            .in3(N__2609),
            .lcout(n13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_idcodeArea_shifter_i9_LC_2_6_3.C_ON=1'b0;
    defparam ctrl_idcodeArea_shifter_i9_LC_2_6_3.SEQ_MODE=4'b1000;
    defparam ctrl_idcodeArea_shifter_i9_LC_2_6_3.LUT_INIT=16'b1111010111011101;
    LogicCell40 ctrl_idcodeArea_shifter_i9_LC_2_6_3 (
            .in0(N__4897),
            .in1(N__3066),
            .in2(N__2598),
            .in3(N__5063),
            .lcout(ctrl_idcodeArea_shifter_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4700),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_idcodeArea_shifter_i11_LC_2_6_4.C_ON=1'b0;
    defparam ctrl_idcodeArea_shifter_i11_LC_2_6_4.SEQ_MODE=4'b1000;
    defparam ctrl_idcodeArea_shifter_i11_LC_2_6_4.LUT_INIT=16'b1101100000000000;
    LogicCell40 ctrl_idcodeArea_shifter_i11_LC_2_6_4 (
            .in0(N__5061),
            .in1(N__3074),
            .in2(N__5112),
            .in3(N__4898),
            .lcout(ctrl_idcodeArea_shifter_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4700),
            .ce(),
            .sr(_gnd_net_));
    defparam i3_2_lut_LC_2_6_6.C_ON=1'b0;
    defparam i3_2_lut_LC_2_6_6.SEQ_MODE=4'b0000;
    defparam i3_2_lut_LC_2_6_6.LUT_INIT=16'b1111111111001100;
    LogicCell40 i3_2_lut_LC_2_6_6 (
            .in0(_gnd_net_),
            .in1(N__2582),
            .in2(_gnd_net_),
            .in3(N__2571),
            .lcout(n11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_idcodeArea_shifter_i10_LC_2_6_7.C_ON=1'b0;
    defparam ctrl_idcodeArea_shifter_i10_LC_2_6_7.SEQ_MODE=4'b1000;
    defparam ctrl_idcodeArea_shifter_i10_LC_2_6_7.LUT_INIT=16'b1000100010100000;
    LogicCell40 ctrl_idcodeArea_shifter_i10_LC_2_6_7 (
            .in0(N__4896),
            .in1(N__3065),
            .in2(N__3078),
            .in3(N__5062),
            .lcout(ctrl_idcodeArea_shifter_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4700),
            .ce(),
            .sr(_gnd_net_));
    defparam i1373_4_lut_LC_2_7_0.C_ON=1'b0;
    defparam i1373_4_lut_LC_2_7_0.SEQ_MODE=4'b0000;
    defparam i1373_4_lut_LC_2_7_0.LUT_INIT=16'b1000000000000000;
    LogicCell40 i1373_4_lut_LC_2_7_0 (
            .in0(N__3056),
            .in1(N__3044),
            .in2(N__3033),
            .in3(N__3017),
            .lcout(n2176),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1357_4_lut_LC_2_7_1.C_ON=1'b0;
    defparam i1357_4_lut_LC_2_7_1.SEQ_MODE=4'b0000;
    defparam i1357_4_lut_LC_2_7_1.LUT_INIT=16'b1000000000000000;
    LogicCell40 i1357_4_lut_LC_2_7_1 (
            .in0(N__3005),
            .in1(N__2993),
            .in2(N__2982),
            .in3(N__2966),
            .lcout(),
            .ltout(n2160_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1379_4_lut_LC_2_7_2.C_ON=1'b0;
    defparam i1379_4_lut_LC_2_7_2.SEQ_MODE=4'b0000;
    defparam i1379_4_lut_LC_2_7_2.LUT_INIT=16'b1000000000000000;
    LogicCell40 i1379_4_lut_LC_2_7_2 (
            .in0(N__2955),
            .in1(N__2766),
            .in2(N__2949),
            .in3(N__2946),
            .lcout(),
            .ltout(n2182_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i7_4_lut_LC_2_7_3.C_ON=1'b0;
    defparam i7_4_lut_LC_2_7_3.SEQ_MODE=4'b0000;
    defparam i7_4_lut_LC_2_7_3.LUT_INIT=16'b1111111111101111;
    LogicCell40 i7_4_lut_LC_2_7_3 (
            .in0(N__2939),
            .in1(N__2928),
            .in2(N__2922),
            .in3(N__2919),
            .lcout(n2113),
            .ltout(n2113_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i990_2_lut_LC_2_7_4.C_ON=1'b0;
    defparam i990_2_lut_LC_2_7_4.SEQ_MODE=4'b0000;
    defparam i990_2_lut_LC_2_7_4.LUT_INIT=16'b0000000011110000;
    LogicCell40 i990_2_lut_LC_2_7_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__2913),
            .in3(N__5261),
            .lcout(n1771),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1359_4_lut_LC_2_7_5.C_ON=1'b0;
    defparam i1359_4_lut_LC_2_7_5.SEQ_MODE=4'b0000;
    defparam i1359_4_lut_LC_2_7_5.LUT_INIT=16'b1000000000000000;
    LogicCell40 i1359_4_lut_LC_2_7_5 (
            .in0(N__2816),
            .in1(N__2804),
            .in2(N__2793),
            .in3(N__2777),
            .lcout(n2162),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam myClockArea_timeout_state_88_LC_2_8_0.C_ON=1'b0;
    defparam myClockArea_timeout_state_88_LC_2_8_0.SEQ_MODE=4'b1010;
    defparam myClockArea_timeout_state_88_LC_2_8_0.LUT_INIT=16'b0000000000110011;
    LogicCell40 myClockArea_timeout_state_88_LC_2_8_0 (
            .in0(_gnd_net_),
            .in1(N__5257),
            .in2(_gnd_net_),
            .in3(N__2760),
            .lcout(myClockArea_timeout_state),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5214),
            .ce(),
            .sr(N__3485));
    defparam ctrl_tap_instructionShift_i0_i1_LC_4_1_0.C_ON=1'b0;
    defparam ctrl_tap_instructionShift_i0_i1_LC_4_1_0.SEQ_MODE=4'b1000;
    defparam ctrl_tap_instructionShift_i0_i1_LC_4_1_0.LUT_INIT=16'b1110111001000100;
    LogicCell40 ctrl_tap_instructionShift_i0_i1_LC_4_1_0 (
            .in0(N__4217),
            .in1(N__3371),
            .in2(_gnd_net_),
            .in3(N__3435),
            .lcout(ctrl_tap_instructionShift_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4714),
            .ce(N__3594),
            .sr(_gnd_net_));
    defparam ctrl_tap_instructionShift_i0_i2_LC_4_1_1.C_ON=1'b0;
    defparam ctrl_tap_instructionShift_i0_i2_LC_4_1_1.SEQ_MODE=4'b1000;
    defparam ctrl_tap_instructionShift_i0_i2_LC_4_1_1.LUT_INIT=16'b1100110010101010;
    LogicCell40 ctrl_tap_instructionShift_i0_i2_LC_4_1_1 (
            .in0(N__3218),
            .in1(N__3404),
            .in2(_gnd_net_),
            .in3(N__4222),
            .lcout(ctrl_tap_instructionShift_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4714),
            .ce(N__3594),
            .sr(_gnd_net_));
    defparam ctrl_tap_instructionShift_i0_i4_LC_4_1_2.C_ON=1'b0;
    defparam ctrl_tap_instructionShift_i0_i4_LC_4_1_2.SEQ_MODE=4'b1000;
    defparam ctrl_tap_instructionShift_i0_i4_LC_4_1_2.LUT_INIT=16'b1110111001000100;
    LogicCell40 ctrl_tap_instructionShift_i0_i4_LC_4_1_2 (
            .in0(N__4218),
            .in1(N__3311),
            .in2(_gnd_net_),
            .in3(N__3359),
            .lcout(ctrl_tap_instructionShift_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4714),
            .ce(N__3594),
            .sr(_gnd_net_));
    defparam ctrl_tap_instructionShift_i0_i5_LC_4_1_3.C_ON=1'b0;
    defparam ctrl_tap_instructionShift_i0_i5_LC_4_1_3.SEQ_MODE=4'b1000;
    defparam ctrl_tap_instructionShift_i0_i5_LC_4_1_3.LUT_INIT=16'b1110111000100010;
    LogicCell40 ctrl_tap_instructionShift_i0_i5_LC_4_1_3 (
            .in0(N__3164),
            .in1(N__4221),
            .in2(_gnd_net_),
            .in3(N__3339),
            .lcout(ctrl_tap_instructionShift_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4714),
            .ce(N__3594),
            .sr(_gnd_net_));
    defparam ctrl_tap_instructionShift_i0_i7_LC_4_1_4.C_ON=1'b0;
    defparam ctrl_tap_instructionShift_i0_i7_LC_4_1_4.SEQ_MODE=4'b1000;
    defparam ctrl_tap_instructionShift_i0_i7_LC_4_1_4.LUT_INIT=16'b1110111001000100;
    LogicCell40 ctrl_tap_instructionShift_i0_i7_LC_4_1_4 (
            .in0(N__4220),
            .in1(N__5181),
            .in2(_gnd_net_),
            .in3(N__3299),
            .lcout(ctrl_tap_instructionShift_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4714),
            .ce(N__3594),
            .sr(_gnd_net_));
    defparam ctrl_tap_instructionShift_i0_i3_LC_4_1_5.C_ON=1'b0;
    defparam ctrl_tap_instructionShift_i0_i3_LC_4_1_5.SEQ_MODE=4'b1000;
    defparam ctrl_tap_instructionShift_i0_i3_LC_4_1_5.LUT_INIT=16'b1100110010101010;
    LogicCell40 ctrl_tap_instructionShift_i0_i3_LC_4_1_5 (
            .in0(N__3263),
            .in1(N__3252),
            .in2(_gnd_net_),
            .in3(N__4223),
            .lcout(ctrl_tap_instructionShift_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4714),
            .ce(N__3594),
            .sr(_gnd_net_));
    defparam ctrl_tap_instructionShift_i0_i6_LC_4_1_6.C_ON=1'b0;
    defparam ctrl_tap_instructionShift_i0_i6_LC_4_1_6.SEQ_MODE=4'b1000;
    defparam ctrl_tap_instructionShift_i0_i6_LC_4_1_6.LUT_INIT=16'b1110111001000100;
    LogicCell40 ctrl_tap_instructionShift_i0_i6_LC_4_1_6 (
            .in0(N__4219),
            .in1(N__3203),
            .in2(_gnd_net_),
            .in3(N__3192),
            .lcout(ctrl_tap_instructionShift_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4714),
            .ce(N__3594),
            .sr(_gnd_net_));
    defparam ctrl_tap_instructionShift_i0_i0_LC_4_2_1.C_ON=1'b0;
    defparam ctrl_tap_instructionShift_i0_i0_LC_4_2_1.SEQ_MODE=4'b1000;
    defparam ctrl_tap_instructionShift_i0_i0_LC_4_2_1.LUT_INIT=16'b1100110010101010;
    LogicCell40 ctrl_tap_instructionShift_i0_i0_LC_4_2_1 (
            .in0(N__3146),
            .in1(N__3135),
            .in2(_gnd_net_),
            .in3(N__4224),
            .lcout(ctrl_tap_instructionShift_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4712),
            .ce(N__3590),
            .sr(_gnd_net_));
    defparam i1436_2_lut_3_lut_4_lut_LC_4_3_0.C_ON=1'b0;
    defparam i1436_2_lut_3_lut_4_lut_LC_4_3_0.SEQ_MODE=4'b0000;
    defparam i1436_2_lut_3_lut_4_lut_LC_4_3_0.LUT_INIT=16'b0000001000000000;
    LogicCell40 i1436_2_lut_3_lut_4_lut_LC_4_3_0 (
            .in0(N__4086),
            .in1(N__3768),
            .in2(N__3702),
            .in3(N__3881),
            .lcout(n1353),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_idcodeArea_shifter_i18_LC_4_3_1.C_ON=1'b0;
    defparam ctrl_idcodeArea_shifter_i18_LC_4_3_1.SEQ_MODE=4'b1000;
    defparam ctrl_idcodeArea_shifter_i18_LC_4_3_1.LUT_INIT=16'b1101111110001111;
    LogicCell40 ctrl_idcodeArea_shifter_i18_LC_4_3_1 (
            .in0(N__5049),
            .in1(N__3746),
            .in2(N__4928),
            .in3(N__3726),
            .lcout(ctrl_idcodeArea_shifter_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4711),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_idcodeArea_shifter_i17_LC_4_3_2.C_ON=1'b0;
    defparam ctrl_idcodeArea_shifter_i17_LC_4_3_2.SEQ_MODE=4'b1000;
    defparam ctrl_idcodeArea_shifter_i17_LC_4_3_2.LUT_INIT=16'b1000100011000000;
    LogicCell40 ctrl_idcodeArea_shifter_i17_LC_4_3_2 (
            .in0(N__5144),
            .in1(N__4900),
            .in2(N__3750),
            .in3(N__5053),
            .lcout(ctrl_idcodeArea_shifter_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4711),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_idcodeArea_shifter_i20_LC_4_3_3.C_ON=1'b0;
    defparam ctrl_idcodeArea_shifter_i20_LC_4_3_3.SEQ_MODE=4'b1000;
    defparam ctrl_idcodeArea_shifter_i20_LC_4_3_3.LUT_INIT=16'b1110010000000000;
    LogicCell40 ctrl_idcodeArea_shifter_i20_LC_4_3_3 (
            .in0(N__5050),
            .in1(N__3555),
            .in2(N__3738),
            .in3(N__4911),
            .lcout(ctrl_idcodeArea_shifter_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4711),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_idcodeArea_shifter_i19_LC_4_3_4.C_ON=1'b0;
    defparam ctrl_idcodeArea_shifter_i19_LC_4_3_4.SEQ_MODE=4'b1000;
    defparam ctrl_idcodeArea_shifter_i19_LC_4_3_4.LUT_INIT=16'b1010110000000000;
    LogicCell40 ctrl_idcodeArea_shifter_i19_LC_4_3_4 (
            .in0(N__3725),
            .in1(N__3737),
            .in2(N__5077),
            .in3(N__4904),
            .lcout(ctrl_idcodeArea_shifter_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4711),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_idcodeArea_shifter_i31_LC_4_3_5.C_ON=1'b0;
    defparam ctrl_idcodeArea_shifter_i31_LC_4_3_5.SEQ_MODE=4'b1000;
    defparam ctrl_idcodeArea_shifter_i31_LC_4_3_5.LUT_INIT=16'b1101100011111111;
    LogicCell40 ctrl_idcodeArea_shifter_i31_LC_4_3_5 (
            .in0(N__5052),
            .in1(N__3716),
            .in2(N__5195),
            .in3(N__4913),
            .lcout(ctrl_idcodeArea_shifter_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4711),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_4_lut_LC_4_3_6.C_ON=1'b0;
    defparam i1_4_lut_4_lut_LC_4_3_6.SEQ_MODE=4'b0000;
    defparam i1_4_lut_4_lut_LC_4_3_6.LUT_INIT=16'b0000001000010000;
    LogicCell40 i1_4_lut_4_lut_LC_4_3_6 (
            .in0(N__4216),
            .in1(N__4085),
            .in2(N__3701),
            .in3(N__3882),
            .lcout(n1067),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_idcodeArea_shifter_i21_LC_4_3_7.C_ON=1'b0;
    defparam ctrl_idcodeArea_shifter_i21_LC_4_3_7.SEQ_MODE=4'b1000;
    defparam ctrl_idcodeArea_shifter_i21_LC_4_3_7.LUT_INIT=16'b1101100011111111;
    LogicCell40 ctrl_idcodeArea_shifter_i21_LC_4_3_7 (
            .in0(N__5051),
            .in1(N__3554),
            .in2(N__3573),
            .in3(N__4912),
            .lcout(ctrl_idcodeArea_shifter_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4711),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_ledsArea_shifter_i0_i0_LC_4_4_0.C_ON=1'b0;
    defparam ctrl_ledsArea_shifter_i0_i0_LC_4_4_0.SEQ_MODE=4'b1000;
    defparam ctrl_ledsArea_shifter_i0_i0_LC_4_4_0.LUT_INIT=16'b0010001011110000;
    LogicCell40 ctrl_ledsArea_shifter_i0_i0_LC_4_4_0 (
            .in0(N__3539),
            .in1(N__4283),
            .in2(N__4622),
            .in3(N__4365),
            .lcout(ctrl_ledsArea_shifter_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4709),
            .ce(N__4236),
            .sr(_gnd_net_));
    defparam ctrl_ledsArea_shifter_i0_i1_LC_4_4_1.C_ON=1'b0;
    defparam ctrl_ledsArea_shifter_i0_i1_LC_4_4_1.SEQ_MODE=4'b1000;
    defparam ctrl_ledsArea_shifter_i0_i1_LC_4_4_1.LUT_INIT=16'b0100010011100100;
    LogicCell40 ctrl_ledsArea_shifter_i0_i1_LC_4_4_1 (
            .in0(N__4361),
            .in1(N__4571),
            .in2(N__4649),
            .in3(N__4287),
            .lcout(ctrl_ledsArea_shifter_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4709),
            .ce(N__4236),
            .sr(_gnd_net_));
    defparam ctrl_ledsArea_shifter_i0_i2_LC_4_4_2.C_ON=1'b0;
    defparam ctrl_ledsArea_shifter_i0_i2_LC_4_4_2.SEQ_MODE=4'b1000;
    defparam ctrl_ledsArea_shifter_i0_i2_LC_4_4_2.LUT_INIT=16'b0010001011110000;
    LogicCell40 ctrl_ledsArea_shifter_i0_i2_LC_4_4_2 (
            .in0(N__4595),
            .in1(N__4284),
            .in2(N__4520),
            .in3(N__4366),
            .lcout(ctrl_ledsArea_shifter_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4709),
            .ce(N__4236),
            .sr(_gnd_net_));
    defparam ctrl_ledsArea_shifter_i0_i3_LC_4_4_3.C_ON=1'b0;
    defparam ctrl_ledsArea_shifter_i0_i3_LC_4_4_3.SEQ_MODE=4'b1000;
    defparam ctrl_ledsArea_shifter_i0_i3_LC_4_4_3.LUT_INIT=16'b0101000011011000;
    LogicCell40 ctrl_ledsArea_shifter_i0_i3_LC_4_4_3 (
            .in0(N__4362),
            .in1(N__4544),
            .in2(N__4481),
            .in3(N__4288),
            .lcout(ctrl_ledsArea_shifter_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4709),
            .ce(N__4236),
            .sr(_gnd_net_));
    defparam ctrl_ledsArea_shifter_i0_i4_LC_4_4_4.C_ON=1'b0;
    defparam ctrl_ledsArea_shifter_i0_i4_LC_4_4_4.SEQ_MODE=4'b1000;
    defparam ctrl_ledsArea_shifter_i0_i4_LC_4_4_4.LUT_INIT=16'b0010111100100000;
    LogicCell40 ctrl_ledsArea_shifter_i0_i4_LC_4_4_4 (
            .in0(N__4503),
            .in1(N__4285),
            .in2(N__4371),
            .in3(N__4427),
            .lcout(ctrl_ledsArea_shifter_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4709),
            .ce(N__4236),
            .sr(_gnd_net_));
    defparam ctrl_ledsArea_shifter_i0_i5_LC_4_4_5.C_ON=1'b0;
    defparam ctrl_ledsArea_shifter_i0_i5_LC_4_4_5.SEQ_MODE=4'b1000;
    defparam ctrl_ledsArea_shifter_i0_i5_LC_4_4_5.LUT_INIT=16'b0101000011011000;
    LogicCell40 ctrl_ledsArea_shifter_i0_i5_LC_4_4_5 (
            .in0(N__4363),
            .in1(N__4457),
            .in2(N__4388),
            .in3(N__4289),
            .lcout(ctrl_ledsArea_shifter_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4709),
            .ce(N__4236),
            .sr(_gnd_net_));
    defparam ctrl_ledsArea_shifter_i0_i6_LC_4_4_6.C_ON=1'b0;
    defparam ctrl_ledsArea_shifter_i0_i6_LC_4_4_6.SEQ_MODE=4'b1000;
    defparam ctrl_ledsArea_shifter_i0_i6_LC_4_4_6.LUT_INIT=16'b0010001011110000;
    LogicCell40 ctrl_ledsArea_shifter_i0_i6_LC_4_4_6 (
            .in0(N__4416),
            .in1(N__4286),
            .in2(N__4253),
            .in3(N__4367),
            .lcout(ctrl_ledsArea_shifter_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4709),
            .ce(N__4236),
            .sr(_gnd_net_));
    defparam ctrl_ledsArea_shifter_i0_i7_LC_4_4_7.C_ON=1'b0;
    defparam ctrl_ledsArea_shifter_i0_i7_LC_4_4_7.SEQ_MODE=4'b1000;
    defparam ctrl_ledsArea_shifter_i0_i7_LC_4_4_7.LUT_INIT=16'b0101000011011000;
    LogicCell40 ctrl_ledsArea_shifter_i0_i7_LC_4_4_7 (
            .in0(N__4364),
            .in1(N__4313),
            .in2(N__5196),
            .in3(N__4290),
            .lcout(ctrl_ledsArea_shifter_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4709),
            .ce(N__4236),
            .sr(_gnd_net_));
    defparam mux_210_i3_4_lut_4_lut_LC_4_5_2.C_ON=1'b0;
    defparam mux_210_i3_4_lut_4_lut_LC_4_5_2.SEQ_MODE=4'b0000;
    defparam mux_210_i3_4_lut_4_lut_LC_4_5_2.LUT_INIT=16'b1101001100010011;
    LogicCell40 mux_210_i3_4_lut_4_lut_LC_4_5_2 (
            .in0(N__4215),
            .in1(N__4084),
            .in2(N__3933),
            .in3(N__3880),
            .lcout(n963),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam myClockArea_toggle_90_LC_4_8_5.C_ON=1'b0;
    defparam myClockArea_toggle_90_LC_4_8_5.SEQ_MODE=4'b1000;
    defparam myClockArea_toggle_90_LC_4_8_5.LUT_INIT=16'b0011001111001100;
    LogicCell40 myClockArea_toggle_90_LC_4_8_5 (
            .in0(_gnd_net_),
            .in1(N__5228),
            .in2(_gnd_net_),
            .in3(N__5262),
            .lcout(io_leds_c_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5217),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_tap_bypass_81_LC_5_2_7.C_ON=1'b0;
    defparam ctrl_tap_bypass_81_LC_5_2_7.SEQ_MODE=4'b1000;
    defparam ctrl_tap_bypass_81_LC_5_2_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 ctrl_tap_bypass_81_LC_5_2_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5185),
            .lcout(ctrl_tap_bypass),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4715),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_idcodeArea_shifter_i14_LC_5_3_0.C_ON=1'b0;
    defparam ctrl_idcodeArea_shifter_i14_LC_5_3_0.SEQ_MODE=4'b1000;
    defparam ctrl_idcodeArea_shifter_i14_LC_5_3_0.LUT_INIT=16'b1101100011111111;
    LogicCell40 ctrl_idcodeArea_shifter_i14_LC_5_3_0 (
            .in0(N__5055),
            .in1(N__5132),
            .in2(N__4728),
            .in3(N__4914),
            .lcout(ctrl_idcodeArea_shifter_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4713),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_idcodeArea_shifter_i16_LC_5_3_1.C_ON=1'b0;
    defparam ctrl_idcodeArea_shifter_i16_LC_5_3_1.SEQ_MODE=4'b1000;
    defparam ctrl_idcodeArea_shifter_i16_LC_5_3_1.LUT_INIT=16'b1011101111110011;
    LogicCell40 ctrl_idcodeArea_shifter_i16_LC_5_3_1 (
            .in0(N__5090),
            .in1(N__4906),
            .in2(N__5148),
            .in3(N__5057),
            .lcout(ctrl_idcodeArea_shifter_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4713),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_idcodeArea_shifter_i13_LC_5_3_2.C_ON=1'b0;
    defparam ctrl_idcodeArea_shifter_i13_LC_5_3_2.SEQ_MODE=4'b1000;
    defparam ctrl_idcodeArea_shifter_i13_LC_5_3_2.LUT_INIT=16'b1101000010000000;
    LogicCell40 ctrl_idcodeArea_shifter_i13_LC_5_3_2 (
            .in0(N__5054),
            .in1(N__5120),
            .in2(N__4929),
            .in3(N__5133),
            .lcout(ctrl_idcodeArea_shifter_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4713),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_idcodeArea_shifter_i12_LC_5_3_3.C_ON=1'b0;
    defparam ctrl_idcodeArea_shifter_i12_LC_5_3_3.SEQ_MODE=4'b1000;
    defparam ctrl_idcodeArea_shifter_i12_LC_5_3_3.LUT_INIT=16'b1000100011000000;
    LogicCell40 ctrl_idcodeArea_shifter_i12_LC_5_3_3 (
            .in0(N__5102),
            .in1(N__4905),
            .in2(N__5124),
            .in3(N__5056),
            .lcout(ctrl_idcodeArea_shifter_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4713),
            .ce(),
            .sr(_gnd_net_));
    defparam ctrl_idcodeArea_shifter_i15_LC_5_3_5.C_ON=1'b0;
    defparam ctrl_idcodeArea_shifter_i15_LC_5_3_5.SEQ_MODE=4'b1000;
    defparam ctrl_idcodeArea_shifter_i15_LC_5_3_5.LUT_INIT=16'b1100101000000000;
    LogicCell40 ctrl_idcodeArea_shifter_i15_LC_5_3_5 (
            .in0(N__5091),
            .in1(N__4727),
            .in2(N__5076),
            .in3(N__4910),
            .lcout(ctrl_idcodeArea_shifter_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4713),
            .ce(),
            .sr(_gnd_net_));
endmodule // MyTopLevel
