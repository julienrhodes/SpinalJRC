-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2017.08.27940

-- Build Date:         Sep 12 2017 08:26:01

-- File Generated:     May 5 2020 16:11:55

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "MyTopLevel" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of MyTopLevel
entity MyTopLevel is
port (
    io_leds : out std_logic_vector(7 downto 0);
    io_jtag_tms : in std_logic;
    io_jtag_tdo : out std_logic;
    io_jtag_tdi : in std_logic;
    io_jtag_tck : in std_logic;
    global_reset : in std_logic;
    global_clk : in std_logic);
end MyTopLevel;

-- Architecture of MyTopLevel
-- View name is \INTERFACE\
architecture \INTERFACE\ of MyTopLevel is

signal \N__4910\ : std_logic;
signal \N__4909\ : std_logic;
signal \N__4908\ : std_logic;
signal \N__4899\ : std_logic;
signal \N__4898\ : std_logic;
signal \N__4897\ : std_logic;
signal \N__4890\ : std_logic;
signal \N__4889\ : std_logic;
signal \N__4888\ : std_logic;
signal \N__4881\ : std_logic;
signal \N__4880\ : std_logic;
signal \N__4879\ : std_logic;
signal \N__4872\ : std_logic;
signal \N__4871\ : std_logic;
signal \N__4870\ : std_logic;
signal \N__4863\ : std_logic;
signal \N__4862\ : std_logic;
signal \N__4861\ : std_logic;
signal \N__4854\ : std_logic;
signal \N__4853\ : std_logic;
signal \N__4852\ : std_logic;
signal \N__4845\ : std_logic;
signal \N__4844\ : std_logic;
signal \N__4843\ : std_logic;
signal \N__4836\ : std_logic;
signal \N__4835\ : std_logic;
signal \N__4834\ : std_logic;
signal \N__4827\ : std_logic;
signal \N__4826\ : std_logic;
signal \N__4825\ : std_logic;
signal \N__4818\ : std_logic;
signal \N__4817\ : std_logic;
signal \N__4816\ : std_logic;
signal \N__4809\ : std_logic;
signal \N__4808\ : std_logic;
signal \N__4807\ : std_logic;
signal \N__4800\ : std_logic;
signal \N__4799\ : std_logic;
signal \N__4798\ : std_logic;
signal \N__4791\ : std_logic;
signal \N__4790\ : std_logic;
signal \N__4789\ : std_logic;
signal \N__4772\ : std_logic;
signal \N__4769\ : std_logic;
signal \N__4766\ : std_logic;
signal \N__4763\ : std_logic;
signal \N__4762\ : std_logic;
signal \N__4759\ : std_logic;
signal \N__4756\ : std_logic;
signal \N__4755\ : std_logic;
signal \N__4752\ : std_logic;
signal \N__4749\ : std_logic;
signal \N__4746\ : std_logic;
signal \N__4739\ : std_logic;
signal \N__4738\ : std_logic;
signal \N__4735\ : std_logic;
signal \N__4732\ : std_logic;
signal \N__4729\ : std_logic;
signal \N__4724\ : std_logic;
signal \N__4721\ : std_logic;
signal \N__4720\ : std_logic;
signal \N__4717\ : std_logic;
signal \N__4714\ : std_logic;
signal \N__4709\ : std_logic;
signal \N__4708\ : std_logic;
signal \N__4705\ : std_logic;
signal \N__4702\ : std_logic;
signal \N__4697\ : std_logic;
signal \N__4696\ : std_logic;
signal \N__4693\ : std_logic;
signal \N__4690\ : std_logic;
signal \N__4687\ : std_logic;
signal \N__4684\ : std_logic;
signal \N__4681\ : std_logic;
signal \N__4678\ : std_logic;
signal \N__4677\ : std_logic;
signal \N__4672\ : std_logic;
signal \N__4669\ : std_logic;
signal \N__4664\ : std_logic;
signal \N__4663\ : std_logic;
signal \N__4660\ : std_logic;
signal \N__4657\ : std_logic;
signal \N__4654\ : std_logic;
signal \N__4651\ : std_logic;
signal \N__4648\ : std_logic;
signal \N__4643\ : std_logic;
signal \N__4642\ : std_logic;
signal \N__4639\ : std_logic;
signal \N__4636\ : std_logic;
signal \N__4633\ : std_logic;
signal \N__4628\ : std_logic;
signal \N__4627\ : std_logic;
signal \N__4626\ : std_logic;
signal \N__4625\ : std_logic;
signal \N__4624\ : std_logic;
signal \N__4619\ : std_logic;
signal \N__4612\ : std_logic;
signal \N__4607\ : std_logic;
signal \N__4604\ : std_logic;
signal \N__4601\ : std_logic;
signal \N__4600\ : std_logic;
signal \N__4597\ : std_logic;
signal \N__4594\ : std_logic;
signal \N__4591\ : std_logic;
signal \N__4588\ : std_logic;
signal \N__4583\ : std_logic;
signal \N__4582\ : std_logic;
signal \N__4579\ : std_logic;
signal \N__4576\ : std_logic;
signal \N__4571\ : std_logic;
signal \N__4570\ : std_logic;
signal \N__4567\ : std_logic;
signal \N__4564\ : std_logic;
signal \N__4561\ : std_logic;
signal \N__4558\ : std_logic;
signal \N__4557\ : std_logic;
signal \N__4556\ : std_logic;
signal \N__4555\ : std_logic;
signal \N__4554\ : std_logic;
signal \N__4553\ : std_logic;
signal \N__4552\ : std_logic;
signal \N__4551\ : std_logic;
signal \N__4548\ : std_logic;
signal \N__4545\ : std_logic;
signal \N__4534\ : std_logic;
signal \N__4529\ : std_logic;
signal \N__4520\ : std_logic;
signal \N__4517\ : std_logic;
signal \N__4514\ : std_logic;
signal \N__4513\ : std_logic;
signal \N__4510\ : std_logic;
signal \N__4507\ : std_logic;
signal \N__4502\ : std_logic;
signal \N__4499\ : std_logic;
signal \N__4498\ : std_logic;
signal \N__4497\ : std_logic;
signal \N__4494\ : std_logic;
signal \N__4491\ : std_logic;
signal \N__4488\ : std_logic;
signal \N__4485\ : std_logic;
signal \N__4482\ : std_logic;
signal \N__4479\ : std_logic;
signal \N__4472\ : std_logic;
signal \N__4471\ : std_logic;
signal \N__4468\ : std_logic;
signal \N__4465\ : std_logic;
signal \N__4462\ : std_logic;
signal \N__4457\ : std_logic;
signal \N__4454\ : std_logic;
signal \N__4451\ : std_logic;
signal \N__4450\ : std_logic;
signal \N__4449\ : std_logic;
signal \N__4446\ : std_logic;
signal \N__4443\ : std_logic;
signal \N__4440\ : std_logic;
signal \N__4433\ : std_logic;
signal \N__4430\ : std_logic;
signal \N__4429\ : std_logic;
signal \N__4426\ : std_logic;
signal \N__4423\ : std_logic;
signal \N__4418\ : std_logic;
signal \N__4417\ : std_logic;
signal \N__4416\ : std_logic;
signal \N__4415\ : std_logic;
signal \N__4414\ : std_logic;
signal \N__4411\ : std_logic;
signal \N__4408\ : std_logic;
signal \N__4405\ : std_logic;
signal \N__4402\ : std_logic;
signal \N__4401\ : std_logic;
signal \N__4400\ : std_logic;
signal \N__4397\ : std_logic;
signal \N__4394\ : std_logic;
signal \N__4393\ : std_logic;
signal \N__4388\ : std_logic;
signal \N__4385\ : std_logic;
signal \N__4380\ : std_logic;
signal \N__4377\ : std_logic;
signal \N__4374\ : std_logic;
signal \N__4371\ : std_logic;
signal \N__4364\ : std_logic;
signal \N__4355\ : std_logic;
signal \N__4352\ : std_logic;
signal \N__4351\ : std_logic;
signal \N__4348\ : std_logic;
signal \N__4345\ : std_logic;
signal \N__4342\ : std_logic;
signal \N__4339\ : std_logic;
signal \N__4338\ : std_logic;
signal \N__4335\ : std_logic;
signal \N__4332\ : std_logic;
signal \N__4329\ : std_logic;
signal \N__4322\ : std_logic;
signal \N__4321\ : std_logic;
signal \N__4320\ : std_logic;
signal \N__4319\ : std_logic;
signal \N__4318\ : std_logic;
signal \N__4317\ : std_logic;
signal \N__4316\ : std_logic;
signal \N__4315\ : std_logic;
signal \N__4314\ : std_logic;
signal \N__4313\ : std_logic;
signal \N__4312\ : std_logic;
signal \N__4311\ : std_logic;
signal \N__4310\ : std_logic;
signal \N__4309\ : std_logic;
signal \N__4308\ : std_logic;
signal \N__4307\ : std_logic;
signal \N__4306\ : std_logic;
signal \N__4305\ : std_logic;
signal \N__4304\ : std_logic;
signal \N__4265\ : std_logic;
signal \N__4262\ : std_logic;
signal \N__4259\ : std_logic;
signal \N__4258\ : std_logic;
signal \N__4255\ : std_logic;
signal \N__4252\ : std_logic;
signal \N__4247\ : std_logic;
signal \N__4244\ : std_logic;
signal \N__4241\ : std_logic;
signal \N__4238\ : std_logic;
signal \N__4235\ : std_logic;
signal \N__4232\ : std_logic;
signal \N__4231\ : std_logic;
signal \N__4228\ : std_logic;
signal \N__4227\ : std_logic;
signal \N__4226\ : std_logic;
signal \N__4223\ : std_logic;
signal \N__4220\ : std_logic;
signal \N__4215\ : std_logic;
signal \N__4208\ : std_logic;
signal \N__4205\ : std_logic;
signal \N__4204\ : std_logic;
signal \N__4203\ : std_logic;
signal \N__4202\ : std_logic;
signal \N__4201\ : std_logic;
signal \N__4200\ : std_logic;
signal \N__4199\ : std_logic;
signal \N__4198\ : std_logic;
signal \N__4195\ : std_logic;
signal \N__4192\ : std_logic;
signal \N__4189\ : std_logic;
signal \N__4184\ : std_logic;
signal \N__4181\ : std_logic;
signal \N__4178\ : std_logic;
signal \N__4175\ : std_logic;
signal \N__4160\ : std_logic;
signal \N__4157\ : std_logic;
signal \N__4156\ : std_logic;
signal \N__4155\ : std_logic;
signal \N__4154\ : std_logic;
signal \N__4153\ : std_logic;
signal \N__4152\ : std_logic;
signal \N__4145\ : std_logic;
signal \N__4144\ : std_logic;
signal \N__4143\ : std_logic;
signal \N__4142\ : std_logic;
signal \N__4141\ : std_logic;
signal \N__4140\ : std_logic;
signal \N__4137\ : std_logic;
signal \N__4134\ : std_logic;
signal \N__4131\ : std_logic;
signal \N__4128\ : std_logic;
signal \N__4125\ : std_logic;
signal \N__4124\ : std_logic;
signal \N__4123\ : std_logic;
signal \N__4122\ : std_logic;
signal \N__4121\ : std_logic;
signal \N__4120\ : std_logic;
signal \N__4117\ : std_logic;
signal \N__4116\ : std_logic;
signal \N__4115\ : std_logic;
signal \N__4114\ : std_logic;
signal \N__4113\ : std_logic;
signal \N__4112\ : std_logic;
signal \N__4111\ : std_logic;
signal \N__4110\ : std_logic;
signal \N__4107\ : std_logic;
signal \N__4100\ : std_logic;
signal \N__4095\ : std_logic;
signal \N__4092\ : std_logic;
signal \N__4083\ : std_logic;
signal \N__4076\ : std_logic;
signal \N__4067\ : std_logic;
signal \N__4060\ : std_logic;
signal \N__4043\ : std_logic;
signal \N__4042\ : std_logic;
signal \N__4041\ : std_logic;
signal \N__4040\ : std_logic;
signal \N__4039\ : std_logic;
signal \N__4038\ : std_logic;
signal \N__4037\ : std_logic;
signal \N__4036\ : std_logic;
signal \N__4035\ : std_logic;
signal \N__4034\ : std_logic;
signal \N__4033\ : std_logic;
signal \N__4032\ : std_logic;
signal \N__4029\ : std_logic;
signal \N__4028\ : std_logic;
signal \N__4027\ : std_logic;
signal \N__4024\ : std_logic;
signal \N__4023\ : std_logic;
signal \N__4022\ : std_logic;
signal \N__4021\ : std_logic;
signal \N__4018\ : std_logic;
signal \N__4017\ : std_logic;
signal \N__4010\ : std_logic;
signal \N__4007\ : std_logic;
signal \N__4004\ : std_logic;
signal \N__4001\ : std_logic;
signal \N__3996\ : std_logic;
signal \N__3987\ : std_logic;
signal \N__3980\ : std_logic;
signal \N__3973\ : std_logic;
signal \N__3956\ : std_logic;
signal \N__3955\ : std_logic;
signal \N__3954\ : std_logic;
signal \N__3953\ : std_logic;
signal \N__3952\ : std_logic;
signal \N__3951\ : std_logic;
signal \N__3950\ : std_logic;
signal \N__3949\ : std_logic;
signal \N__3946\ : std_logic;
signal \N__3945\ : std_logic;
signal \N__3944\ : std_logic;
signal \N__3943\ : std_logic;
signal \N__3940\ : std_logic;
signal \N__3939\ : std_logic;
signal \N__3934\ : std_logic;
signal \N__3931\ : std_logic;
signal \N__3926\ : std_logic;
signal \N__3923\ : std_logic;
signal \N__3920\ : std_logic;
signal \N__3913\ : std_logic;
signal \N__3912\ : std_logic;
signal \N__3907\ : std_logic;
signal \N__3900\ : std_logic;
signal \N__3897\ : std_logic;
signal \N__3892\ : std_logic;
signal \N__3889\ : std_logic;
signal \N__3886\ : std_logic;
signal \N__3883\ : std_logic;
signal \N__3880\ : std_logic;
signal \N__3877\ : std_logic;
signal \N__3874\ : std_logic;
signal \N__3871\ : std_logic;
signal \N__3868\ : std_logic;
signal \N__3865\ : std_logic;
signal \N__3860\ : std_logic;
signal \N__3851\ : std_logic;
signal \N__3850\ : std_logic;
signal \N__3849\ : std_logic;
signal \N__3848\ : std_logic;
signal \N__3847\ : std_logic;
signal \N__3844\ : std_logic;
signal \N__3843\ : std_logic;
signal \N__3842\ : std_logic;
signal \N__3841\ : std_logic;
signal \N__3840\ : std_logic;
signal \N__3839\ : std_logic;
signal \N__3838\ : std_logic;
signal \N__3837\ : std_logic;
signal \N__3836\ : std_logic;
signal \N__3829\ : std_logic;
signal \N__3826\ : std_logic;
signal \N__3823\ : std_logic;
signal \N__3822\ : std_logic;
signal \N__3821\ : std_logic;
signal \N__3820\ : std_logic;
signal \N__3819\ : std_logic;
signal \N__3818\ : std_logic;
signal \N__3817\ : std_logic;
signal \N__3816\ : std_logic;
signal \N__3815\ : std_logic;
signal \N__3814\ : std_logic;
signal \N__3807\ : std_logic;
signal \N__3804\ : std_logic;
signal \N__3799\ : std_logic;
signal \N__3794\ : std_logic;
signal \N__3791\ : std_logic;
signal \N__3786\ : std_logic;
signal \N__3779\ : std_logic;
signal \N__3774\ : std_logic;
signal \N__3765\ : std_logic;
signal \N__3746\ : std_logic;
signal \N__3743\ : std_logic;
signal \N__3740\ : std_logic;
signal \N__3737\ : std_logic;
signal \N__3734\ : std_logic;
signal \N__3733\ : std_logic;
signal \N__3732\ : std_logic;
signal \N__3731\ : std_logic;
signal \N__3730\ : std_logic;
signal \N__3727\ : std_logic;
signal \N__3726\ : std_logic;
signal \N__3725\ : std_logic;
signal \N__3724\ : std_logic;
signal \N__3723\ : std_logic;
signal \N__3722\ : std_logic;
signal \N__3721\ : std_logic;
signal \N__3720\ : std_logic;
signal \N__3719\ : std_logic;
signal \N__3716\ : std_logic;
signal \N__3715\ : std_logic;
signal \N__3712\ : std_logic;
signal \N__3711\ : std_logic;
signal \N__3708\ : std_logic;
signal \N__3707\ : std_logic;
signal \N__3706\ : std_logic;
signal \N__3705\ : std_logic;
signal \N__3704\ : std_logic;
signal \N__3703\ : std_logic;
signal \N__3700\ : std_logic;
signal \N__3699\ : std_logic;
signal \N__3698\ : std_logic;
signal \N__3697\ : std_logic;
signal \N__3694\ : std_logic;
signal \N__3689\ : std_logic;
signal \N__3680\ : std_logic;
signal \N__3677\ : std_logic;
signal \N__3672\ : std_logic;
signal \N__3669\ : std_logic;
signal \N__3664\ : std_logic;
signal \N__3661\ : std_logic;
signal \N__3656\ : std_logic;
signal \N__3649\ : std_logic;
signal \N__3644\ : std_logic;
signal \N__3639\ : std_logic;
signal \N__3614\ : std_logic;
signal \N__3611\ : std_logic;
signal \N__3608\ : std_logic;
signal \N__3605\ : std_logic;
signal \N__3602\ : std_logic;
signal \N__3599\ : std_logic;
signal \N__3596\ : std_logic;
signal \N__3593\ : std_logic;
signal \N__3590\ : std_logic;
signal \N__3589\ : std_logic;
signal \N__3586\ : std_logic;
signal \N__3583\ : std_logic;
signal \N__3580\ : std_logic;
signal \N__3575\ : std_logic;
signal \N__3572\ : std_logic;
signal \N__3569\ : std_logic;
signal \N__3566\ : std_logic;
signal \N__3563\ : std_logic;
signal \N__3560\ : std_logic;
signal \N__3557\ : std_logic;
signal \N__3554\ : std_logic;
signal \N__3551\ : std_logic;
signal \N__3550\ : std_logic;
signal \N__3547\ : std_logic;
signal \N__3544\ : std_logic;
signal \N__3539\ : std_logic;
signal \N__3538\ : std_logic;
signal \N__3535\ : std_logic;
signal \N__3532\ : std_logic;
signal \N__3527\ : std_logic;
signal \N__3524\ : std_logic;
signal \N__3523\ : std_logic;
signal \N__3522\ : std_logic;
signal \N__3519\ : std_logic;
signal \N__3516\ : std_logic;
signal \N__3513\ : std_logic;
signal \N__3512\ : std_logic;
signal \N__3509\ : std_logic;
signal \N__3506\ : std_logic;
signal \N__3503\ : std_logic;
signal \N__3500\ : std_logic;
signal \N__3495\ : std_logic;
signal \N__3490\ : std_logic;
signal \N__3485\ : std_logic;
signal \N__3484\ : std_logic;
signal \N__3481\ : std_logic;
signal \N__3478\ : std_logic;
signal \N__3475\ : std_logic;
signal \N__3470\ : std_logic;
signal \N__3469\ : std_logic;
signal \N__3466\ : std_logic;
signal \N__3463\ : std_logic;
signal \N__3460\ : std_logic;
signal \N__3455\ : std_logic;
signal \N__3454\ : std_logic;
signal \N__3449\ : std_logic;
signal \N__3446\ : std_logic;
signal \N__3445\ : std_logic;
signal \N__3442\ : std_logic;
signal \N__3439\ : std_logic;
signal \N__3436\ : std_logic;
signal \N__3431\ : std_logic;
signal \N__3430\ : std_logic;
signal \N__3429\ : std_logic;
signal \N__3428\ : std_logic;
signal \N__3427\ : std_logic;
signal \N__3426\ : std_logic;
signal \N__3425\ : std_logic;
signal \N__3424\ : std_logic;
signal \N__3423\ : std_logic;
signal \N__3422\ : std_logic;
signal \N__3421\ : std_logic;
signal \N__3420\ : std_logic;
signal \N__3419\ : std_logic;
signal \N__3418\ : std_logic;
signal \N__3417\ : std_logic;
signal \N__3416\ : std_logic;
signal \N__3415\ : std_logic;
signal \N__3414\ : std_logic;
signal \N__3413\ : std_logic;
signal \N__3412\ : std_logic;
signal \N__3411\ : std_logic;
signal \N__3410\ : std_logic;
signal \N__3409\ : std_logic;
signal \N__3408\ : std_logic;
signal \N__3407\ : std_logic;
signal \N__3406\ : std_logic;
signal \N__3405\ : std_logic;
signal \N__3404\ : std_logic;
signal \N__3403\ : std_logic;
signal \N__3402\ : std_logic;
signal \N__3401\ : std_logic;
signal \N__3400\ : std_logic;
signal \N__3397\ : std_logic;
signal \N__3388\ : std_logic;
signal \N__3371\ : std_logic;
signal \N__3360\ : std_logic;
signal \N__3349\ : std_logic;
signal \N__3332\ : std_logic;
signal \N__3327\ : std_logic;
signal \N__3314\ : std_logic;
signal \N__3313\ : std_logic;
signal \N__3310\ : std_logic;
signal \N__3307\ : std_logic;
signal \N__3302\ : std_logic;
signal \N__3299\ : std_logic;
signal \N__3298\ : std_logic;
signal \N__3297\ : std_logic;
signal \N__3296\ : std_logic;
signal \N__3295\ : std_logic;
signal \N__3294\ : std_logic;
signal \N__3293\ : std_logic;
signal \N__3292\ : std_logic;
signal \N__3291\ : std_logic;
signal \N__3290\ : std_logic;
signal \N__3287\ : std_logic;
signal \N__3286\ : std_logic;
signal \N__3285\ : std_logic;
signal \N__3282\ : std_logic;
signal \N__3279\ : std_logic;
signal \N__3278\ : std_logic;
signal \N__3275\ : std_logic;
signal \N__3272\ : std_logic;
signal \N__3271\ : std_logic;
signal \N__3270\ : std_logic;
signal \N__3267\ : std_logic;
signal \N__3266\ : std_logic;
signal \N__3263\ : std_logic;
signal \N__3260\ : std_logic;
signal \N__3259\ : std_logic;
signal \N__3250\ : std_logic;
signal \N__3249\ : std_logic;
signal \N__3248\ : std_logic;
signal \N__3247\ : std_logic;
signal \N__3246\ : std_logic;
signal \N__3245\ : std_logic;
signal \N__3244\ : std_logic;
signal \N__3243\ : std_logic;
signal \N__3242\ : std_logic;
signal \N__3241\ : std_logic;
signal \N__3240\ : std_logic;
signal \N__3239\ : std_logic;
signal \N__3238\ : std_logic;
signal \N__3237\ : std_logic;
signal \N__3220\ : std_logic;
signal \N__3209\ : std_logic;
signal \N__3208\ : std_logic;
signal \N__3207\ : std_logic;
signal \N__3206\ : std_logic;
signal \N__3205\ : std_logic;
signal \N__3204\ : std_logic;
signal \N__3203\ : std_logic;
signal \N__3200\ : std_logic;
signal \N__3193\ : std_logic;
signal \N__3188\ : std_logic;
signal \N__3179\ : std_logic;
signal \N__3170\ : std_logic;
signal \N__3165\ : std_logic;
signal \N__3160\ : std_logic;
signal \N__3151\ : std_logic;
signal \N__3134\ : std_logic;
signal \N__3133\ : std_logic;
signal \N__3130\ : std_logic;
signal \N__3125\ : std_logic;
signal \N__3122\ : std_logic;
signal \N__3119\ : std_logic;
signal \N__3118\ : std_logic;
signal \N__3117\ : std_logic;
signal \N__3116\ : std_logic;
signal \N__3115\ : std_logic;
signal \N__3114\ : std_logic;
signal \N__3113\ : std_logic;
signal \N__3112\ : std_logic;
signal \N__3111\ : std_logic;
signal \N__3110\ : std_logic;
signal \N__3109\ : std_logic;
signal \N__3108\ : std_logic;
signal \N__3099\ : std_logic;
signal \N__3098\ : std_logic;
signal \N__3097\ : std_logic;
signal \N__3096\ : std_logic;
signal \N__3095\ : std_logic;
signal \N__3094\ : std_logic;
signal \N__3093\ : std_logic;
signal \N__3092\ : std_logic;
signal \N__3091\ : std_logic;
signal \N__3090\ : std_logic;
signal \N__3089\ : std_logic;
signal \N__3088\ : std_logic;
signal \N__3079\ : std_logic;
signal \N__3070\ : std_logic;
signal \N__3067\ : std_logic;
signal \N__3058\ : std_logic;
signal \N__3051\ : std_logic;
signal \N__3042\ : std_logic;
signal \N__3029\ : std_logic;
signal \N__3028\ : std_logic;
signal \N__3025\ : std_logic;
signal \N__3022\ : std_logic;
signal \N__3017\ : std_logic;
signal \N__3016\ : std_logic;
signal \N__3013\ : std_logic;
signal \N__3010\ : std_logic;
signal \N__3005\ : std_logic;
signal \N__3002\ : std_logic;
signal \N__2999\ : std_logic;
signal \N__2998\ : std_logic;
signal \N__2995\ : std_logic;
signal \N__2992\ : std_logic;
signal \N__2987\ : std_logic;
signal \N__2986\ : std_logic;
signal \N__2983\ : std_logic;
signal \N__2980\ : std_logic;
signal \N__2975\ : std_logic;
signal \N__2974\ : std_logic;
signal \N__2971\ : std_logic;
signal \N__2968\ : std_logic;
signal \N__2965\ : std_logic;
signal \N__2960\ : std_logic;
signal \N__2959\ : std_logic;
signal \N__2956\ : std_logic;
signal \N__2953\ : std_logic;
signal \N__2948\ : std_logic;
signal \N__2945\ : std_logic;
signal \N__2942\ : std_logic;
signal \N__2941\ : std_logic;
signal \N__2938\ : std_logic;
signal \N__2935\ : std_logic;
signal \N__2930\ : std_logic;
signal \N__2929\ : std_logic;
signal \N__2926\ : std_logic;
signal \N__2923\ : std_logic;
signal \N__2918\ : std_logic;
signal \N__2917\ : std_logic;
signal \N__2914\ : std_logic;
signal \N__2911\ : std_logic;
signal \N__2908\ : std_logic;
signal \N__2903\ : std_logic;
signal \N__2902\ : std_logic;
signal \N__2899\ : std_logic;
signal \N__2896\ : std_logic;
signal \N__2891\ : std_logic;
signal \N__2888\ : std_logic;
signal \N__2885\ : std_logic;
signal \N__2884\ : std_logic;
signal \N__2883\ : std_logic;
signal \N__2880\ : std_logic;
signal \N__2877\ : std_logic;
signal \N__2874\ : std_logic;
signal \N__2871\ : std_logic;
signal \N__2864\ : std_logic;
signal \N__2861\ : std_logic;
signal \N__2860\ : std_logic;
signal \N__2857\ : std_logic;
signal \N__2854\ : std_logic;
signal \N__2849\ : std_logic;
signal \N__2848\ : std_logic;
signal \N__2847\ : std_logic;
signal \N__2846\ : std_logic;
signal \N__2845\ : std_logic;
signal \N__2834\ : std_logic;
signal \N__2831\ : std_logic;
signal \N__2828\ : std_logic;
signal \N__2827\ : std_logic;
signal \N__2822\ : std_logic;
signal \N__2819\ : std_logic;
signal \N__2818\ : std_logic;
signal \N__2815\ : std_logic;
signal \N__2810\ : std_logic;
signal \N__2807\ : std_logic;
signal \N__2804\ : std_logic;
signal \N__2801\ : std_logic;
signal \N__2800\ : std_logic;
signal \N__2797\ : std_logic;
signal \N__2796\ : std_logic;
signal \N__2793\ : std_logic;
signal \N__2790\ : std_logic;
signal \N__2787\ : std_logic;
signal \N__2784\ : std_logic;
signal \N__2777\ : std_logic;
signal \N__2776\ : std_logic;
signal \N__2773\ : std_logic;
signal \N__2770\ : std_logic;
signal \N__2765\ : std_logic;
signal \N__2764\ : std_logic;
signal \N__2761\ : std_logic;
signal \N__2758\ : std_logic;
signal \N__2753\ : std_logic;
signal \N__2752\ : std_logic;
signal \N__2749\ : std_logic;
signal \N__2746\ : std_logic;
signal \N__2743\ : std_logic;
signal \N__2738\ : std_logic;
signal \N__2737\ : std_logic;
signal \N__2734\ : std_logic;
signal \N__2731\ : std_logic;
signal \N__2726\ : std_logic;
signal \N__2723\ : std_logic;
signal \N__2720\ : std_logic;
signal \N__2719\ : std_logic;
signal \N__2716\ : std_logic;
signal \N__2713\ : std_logic;
signal \N__2708\ : std_logic;
signal \N__2707\ : std_logic;
signal \N__2704\ : std_logic;
signal \N__2701\ : std_logic;
signal \N__2696\ : std_logic;
signal \N__2695\ : std_logic;
signal \N__2692\ : std_logic;
signal \N__2689\ : std_logic;
signal \N__2686\ : std_logic;
signal \N__2681\ : std_logic;
signal \N__2680\ : std_logic;
signal \N__2677\ : std_logic;
signal \N__2674\ : std_logic;
signal \N__2669\ : std_logic;
signal \N__2668\ : std_logic;
signal \N__2665\ : std_logic;
signal \N__2662\ : std_logic;
signal \N__2657\ : std_logic;
signal \N__2656\ : std_logic;
signal \N__2653\ : std_logic;
signal \N__2650\ : std_logic;
signal \N__2645\ : std_logic;
signal \N__2644\ : std_logic;
signal \N__2641\ : std_logic;
signal \N__2638\ : std_logic;
signal \N__2635\ : std_logic;
signal \N__2630\ : std_logic;
signal \N__2629\ : std_logic;
signal \N__2626\ : std_logic;
signal \N__2623\ : std_logic;
signal \N__2618\ : std_logic;
signal \N__2615\ : std_logic;
signal \N__2612\ : std_logic;
signal \N__2609\ : std_logic;
signal \N__2606\ : std_logic;
signal \N__2603\ : std_logic;
signal \N__2602\ : std_logic;
signal \N__2599\ : std_logic;
signal \N__2596\ : std_logic;
signal \N__2591\ : std_logic;
signal \N__2588\ : std_logic;
signal \N__2585\ : std_logic;
signal \N__2582\ : std_logic;
signal \N__2579\ : std_logic;
signal \N__2576\ : std_logic;
signal \N__2573\ : std_logic;
signal \N__2570\ : std_logic;
signal \N__2567\ : std_logic;
signal \N__2566\ : std_logic;
signal \N__2563\ : std_logic;
signal \N__2560\ : std_logic;
signal \N__2557\ : std_logic;
signal \N__2552\ : std_logic;
signal \N__2549\ : std_logic;
signal \N__2546\ : std_logic;
signal \N__2543\ : std_logic;
signal \N__2540\ : std_logic;
signal \N__2537\ : std_logic;
signal \N__2534\ : std_logic;
signal \N__2531\ : std_logic;
signal \N__2528\ : std_logic;
signal \N__2525\ : std_logic;
signal \N__2522\ : std_logic;
signal \N__2521\ : std_logic;
signal \N__2520\ : std_logic;
signal \N__2519\ : std_logic;
signal \N__2518\ : std_logic;
signal \N__2515\ : std_logic;
signal \N__2512\ : std_logic;
signal \N__2509\ : std_logic;
signal \N__2504\ : std_logic;
signal \N__2495\ : std_logic;
signal \N__2492\ : std_logic;
signal \N__2491\ : std_logic;
signal \N__2488\ : std_logic;
signal \N__2485\ : std_logic;
signal \N__2480\ : std_logic;
signal \N__2479\ : std_logic;
signal \N__2476\ : std_logic;
signal \N__2475\ : std_logic;
signal \N__2474\ : std_logic;
signal \N__2471\ : std_logic;
signal \N__2470\ : std_logic;
signal \N__2467\ : std_logic;
signal \N__2464\ : std_logic;
signal \N__2461\ : std_logic;
signal \N__2456\ : std_logic;
signal \N__2447\ : std_logic;
signal \N__2444\ : std_logic;
signal \N__2443\ : std_logic;
signal \N__2440\ : std_logic;
signal \N__2437\ : std_logic;
signal \N__2432\ : std_logic;
signal \N__2431\ : std_logic;
signal \N__2430\ : std_logic;
signal \N__2429\ : std_logic;
signal \N__2428\ : std_logic;
signal \N__2425\ : std_logic;
signal \N__2422\ : std_logic;
signal \N__2419\ : std_logic;
signal \N__2414\ : std_logic;
signal \N__2405\ : std_logic;
signal \N__2404\ : std_logic;
signal \N__2403\ : std_logic;
signal \N__2396\ : std_logic;
signal \N__2393\ : std_logic;
signal \N__2390\ : std_logic;
signal \N__2389\ : std_logic;
signal \N__2386\ : std_logic;
signal \N__2383\ : std_logic;
signal \N__2378\ : std_logic;
signal \N__2377\ : std_logic;
signal \N__2376\ : std_logic;
signal \N__2373\ : std_logic;
signal \N__2372\ : std_logic;
signal \N__2371\ : std_logic;
signal \N__2368\ : std_logic;
signal \N__2365\ : std_logic;
signal \N__2362\ : std_logic;
signal \N__2359\ : std_logic;
signal \N__2356\ : std_logic;
signal \N__2345\ : std_logic;
signal \N__2342\ : std_logic;
signal \N__2339\ : std_logic;
signal \N__2336\ : std_logic;
signal \N__2333\ : std_logic;
signal \N__2332\ : std_logic;
signal \N__2329\ : std_logic;
signal \N__2326\ : std_logic;
signal \N__2323\ : std_logic;
signal \N__2318\ : std_logic;
signal \N__2317\ : std_logic;
signal \N__2314\ : std_logic;
signal \N__2311\ : std_logic;
signal \N__2306\ : std_logic;
signal \N__2303\ : std_logic;
signal \N__2302\ : std_logic;
signal \N__2297\ : std_logic;
signal \N__2294\ : std_logic;
signal \N__2291\ : std_logic;
signal \N__2288\ : std_logic;
signal \N__2285\ : std_logic;
signal \N__2284\ : std_logic;
signal \N__2281\ : std_logic;
signal \N__2278\ : std_logic;
signal \N__2275\ : std_logic;
signal \N__2272\ : std_logic;
signal \N__2267\ : std_logic;
signal \N__2264\ : std_logic;
signal \N__2263\ : std_logic;
signal \N__2260\ : std_logic;
signal \N__2257\ : std_logic;
signal \N__2254\ : std_logic;
signal \N__2249\ : std_logic;
signal \N__2246\ : std_logic;
signal \N__2243\ : std_logic;
signal \N__2240\ : std_logic;
signal \N__2237\ : std_logic;
signal \N__2234\ : std_logic;
signal \N__2231\ : std_logic;
signal \N__2228\ : std_logic;
signal \N__2227\ : std_logic;
signal \N__2224\ : std_logic;
signal \N__2223\ : std_logic;
signal \N__2220\ : std_logic;
signal \N__2217\ : std_logic;
signal \N__2214\ : std_logic;
signal \N__2213\ : std_logic;
signal \N__2210\ : std_logic;
signal \N__2205\ : std_logic;
signal \N__2202\ : std_logic;
signal \N__2195\ : std_logic;
signal \N__2192\ : std_logic;
signal \N__2189\ : std_logic;
signal \N__2186\ : std_logic;
signal \N__2185\ : std_logic;
signal \N__2180\ : std_logic;
signal \N__2177\ : std_logic;
signal \N__2176\ : std_logic;
signal \N__2171\ : std_logic;
signal \N__2168\ : std_logic;
signal \N__2165\ : std_logic;
signal \N__2164\ : std_logic;
signal \N__2159\ : std_logic;
signal \N__2156\ : std_logic;
signal \N__2155\ : std_logic;
signal \N__2150\ : std_logic;
signal \N__2147\ : std_logic;
signal \N__2144\ : std_logic;
signal \N__2141\ : std_logic;
signal \N__2138\ : std_logic;
signal \N__2135\ : std_logic;
signal \N__2132\ : std_logic;
signal \N__2129\ : std_logic;
signal \N__2126\ : std_logic;
signal \N__2123\ : std_logic;
signal \N__2120\ : std_logic;
signal \N__2117\ : std_logic;
signal \N__2114\ : std_logic;
signal \N__2111\ : std_logic;
signal \N__2108\ : std_logic;
signal \N__2105\ : std_logic;
signal \N__2102\ : std_logic;
signal \N__2099\ : std_logic;
signal \N__2096\ : std_logic;
signal \N__2093\ : std_logic;
signal \N__2090\ : std_logic;
signal \N__2087\ : std_logic;
signal \N__2084\ : std_logic;
signal \N__2081\ : std_logic;
signal \N__2078\ : std_logic;
signal \N__2075\ : std_logic;
signal \N__2072\ : std_logic;
signal \N__2069\ : std_logic;
signal \N__2066\ : std_logic;
signal \N__2065\ : std_logic;
signal \N__2060\ : std_logic;
signal \N__2057\ : std_logic;
signal \N__2056\ : std_logic;
signal \N__2053\ : std_logic;
signal \N__2050\ : std_logic;
signal \N__2045\ : std_logic;
signal \N__2042\ : std_logic;
signal \N__2041\ : std_logic;
signal \N__2038\ : std_logic;
signal \N__2033\ : std_logic;
signal \N__2030\ : std_logic;
signal \N__2029\ : std_logic;
signal \N__2026\ : std_logic;
signal \N__2021\ : std_logic;
signal \N__2018\ : std_logic;
signal \N__2017\ : std_logic;
signal \N__2014\ : std_logic;
signal \N__2009\ : std_logic;
signal \N__2006\ : std_logic;
signal \N__2003\ : std_logic;
signal \N__2002\ : std_logic;
signal \N__1999\ : std_logic;
signal \N__1996\ : std_logic;
signal \N__1991\ : std_logic;
signal \N__1990\ : std_logic;
signal \N__1987\ : std_logic;
signal \N__1984\ : std_logic;
signal \N__1979\ : std_logic;
signal \N__1976\ : std_logic;
signal \N__1975\ : std_logic;
signal \N__1970\ : std_logic;
signal \N__1967\ : std_logic;
signal \N__1966\ : std_logic;
signal \N__1963\ : std_logic;
signal \N__1958\ : std_logic;
signal \N__1955\ : std_logic;
signal \N__1954\ : std_logic;
signal \N__1949\ : std_logic;
signal \N__1946\ : std_logic;
signal \N__1945\ : std_logic;
signal \N__1940\ : std_logic;
signal \N__1937\ : std_logic;
signal \N__1936\ : std_logic;
signal \N__1931\ : std_logic;
signal \N__1928\ : std_logic;
signal \N__1925\ : std_logic;
signal \N__1924\ : std_logic;
signal \N__1919\ : std_logic;
signal \N__1916\ : std_logic;
signal \N__1915\ : std_logic;
signal \N__1910\ : std_logic;
signal \N__1907\ : std_logic;
signal \N__1906\ : std_logic;
signal \N__1903\ : std_logic;
signal \N__1900\ : std_logic;
signal \N__1897\ : std_logic;
signal \N__1892\ : std_logic;
signal \N__1889\ : std_logic;
signal \N__1886\ : std_logic;
signal \N__1883\ : std_logic;
signal \N__1880\ : std_logic;
signal \N__1879\ : std_logic;
signal \N__1876\ : std_logic;
signal \N__1873\ : std_logic;
signal \N__1872\ : std_logic;
signal \N__1869\ : std_logic;
signal \N__1866\ : std_logic;
signal \N__1863\ : std_logic;
signal \N__1856\ : std_logic;
signal \N__1853\ : std_logic;
signal \N__1850\ : std_logic;
signal \N__1847\ : std_logic;
signal \N__1844\ : std_logic;
signal \N__1841\ : std_logic;
signal io_jtag_tck_pad_gb_input : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal io_leds_c_0 : std_logic;
signal \ctrl_idcodeArea_shifter_7\ : std_logic;
signal \ctrl_idcodeArea_shifter_10\ : std_logic;
signal \ctrl_idcodeArea_shifter_9\ : std_logic;
signal \ctrl_idcodeArea_shifter_8\ : std_logic;
signal \ctrl_idcodeArea_shifter_4\ : std_logic;
signal \ctrl_idcodeArea_shifter_6\ : std_logic;
signal \ctrl_idcodeArea_shifter_5\ : std_logic;
signal \ctrl_idcodeArea_shifter_11\ : std_logic;
signal \ctrl_idcodeArea_shifter_16\ : std_logic;
signal \ctrl_idcodeArea_shifter_15\ : std_logic;
signal \ctrl_idcodeArea_shifter_14\ : std_logic;
signal \ctrl_idcodeArea_shifter_13\ : std_logic;
signal \ctrl_idcodeArea_shifter_12\ : std_logic;
signal \ctrl_idcodeArea_shifter_3\ : std_logic;
signal \ctrl_idcodeArea_shifter_2\ : std_logic;
signal n7 : std_logic;
signal \n7_cascade_\ : std_logic;
signal n2206 : std_logic;
signal \n7_adj_1_cascade_\ : std_logic;
signal \bfn_4_7_0_\ : std_logic;
signal n2059 : std_logic;
signal n2060 : std_logic;
signal n2061 : std_logic;
signal n2062 : std_logic;
signal n2063 : std_logic;
signal n2064 : std_logic;
signal n2065 : std_logic;
signal n2066 : std_logic;
signal \bfn_4_8_0_\ : std_logic;
signal n2067 : std_logic;
signal n2068 : std_logic;
signal n2069 : std_logic;
signal n2070 : std_logic;
signal n2071 : std_logic;
signal n2072 : std_logic;
signal n2073 : std_logic;
signal n2074 : std_logic;
signal \bfn_4_9_0_\ : std_logic;
signal n2075 : std_logic;
signal n2076 : std_logic;
signal n2077 : std_logic;
signal n2078 : std_logic;
signal n2079 : std_logic;
signal n2080 : std_logic;
signal global_reset_c : std_logic;
signal \ctrl_idcodeArea_shifter_31\ : std_logic;
signal \ctrl_idcodeArea_shifter_28\ : std_logic;
signal \ctrl_idcodeArea_shifter_30\ : std_logic;
signal \ctrl_idcodeArea_shifter_29\ : std_logic;
signal \ctrl_idcodeArea_shifter_17\ : std_logic;
signal \ctrl_idcodeArea_shifter_1\ : std_logic;
signal \n6_cascade_\ : std_logic;
signal \ctrl_idcodeArea_shifter_0\ : std_logic;
signal n2085 : std_logic;
signal \n15_cascade_\ : std_logic;
signal n7_adj_1 : std_logic;
signal \ctrl_ledsArea_shifter_0\ : std_logic;
signal \ctrl_tap_tdoUnbufferd_N_211_cascade_\ : std_logic;
signal \ctrl_tap_tdoUnbufferd\ : std_logic;
signal \n1489_cascade_\ : std_logic;
signal \n1269_cascade_\ : std_logic;
signal ctrl_tap_instruction_0 : std_logic;
signal \ctrl_tap_instructionShift_3\ : std_logic;
signal ctrl_tap_instruction_3 : std_logic;
signal \ctrl_tap_instructionShift_2\ : std_logic;
signal ctrl_tap_instruction_2 : std_logic;
signal n1269 : std_logic;
signal \ctrl_tap_instructionShift_1\ : std_logic;
signal ctrl_tap_instruction_1 : std_logic;
signal n2248 : std_logic;
signal \n118_cascade_\ : std_logic;
signal \n2282_cascade_\ : std_logic;
signal \n2326_cascade_\ : std_logic;
signal n2306 : std_logic;
signal n1022 : std_logic;
signal \n2231_cascade_\ : std_logic;
signal n2273 : std_logic;
signal \n2263_cascade_\ : std_logic;
signal n2323 : std_logic;
signal n2272 : std_logic;
signal io_leds_c_7 : std_logic;
signal \myClockArea_timeout_counter_value_3\ : std_logic;
signal \myClockArea_timeout_counter_value_1\ : std_logic;
signal \myClockArea_timeout_counter_value_5\ : std_logic;
signal \myClockArea_timeout_counter_value_0\ : std_logic;
signal n2309 : std_logic;
signal \myClockArea_timeout_counter_value_4\ : std_logic;
signal \myClockArea_timeout_counter_value_6\ : std_logic;
signal \myClockArea_timeout_counter_value_22\ : std_logic;
signal \myClockArea_timeout_counter_value_16\ : std_logic;
signal \myClockArea_timeout_counter_value_17\ : std_logic;
signal \myClockArea_timeout_counter_value_8\ : std_logic;
signal \myClockArea_timeout_counter_value_10\ : std_logic;
signal \myClockArea_timeout_counter_value_2\ : std_logic;
signal n2216 : std_logic;
signal \n2218_cascade_\ : std_logic;
signal n2222 : std_logic;
signal \myClockArea_timeout_counter_value_13\ : std_logic;
signal \n2228_cascade_\ : std_logic;
signal n2185 : std_logic;
signal \n2185_cascade_\ : std_logic;
signal n1848 : std_logic;
signal \myClockArea_timeout_counter_value_7\ : std_logic;
signal \myClockArea_timeout_counter_value_21\ : std_logic;
signal n11 : std_logic;
signal \myClockArea_timeout_counter_value_19\ : std_logic;
signal \myClockArea_timeout_counter_value_15\ : std_logic;
signal \myClockArea_timeout_counter_value_20\ : std_logic;
signal \myClockArea_timeout_counter_value_11\ : std_logic;
signal n2220 : std_logic;
signal \myClockArea_timeout_counter_value_9\ : std_logic;
signal \myClockArea_timeout_counter_value_18\ : std_logic;
signal \myClockArea_timeout_counter_value_12\ : std_logic;
signal \myClockArea_timeout_counter_value_14\ : std_logic;
signal n13 : std_logic;
signal \myClockArea_timeout_state\ : std_logic;
signal io_leds_c_3 : std_logic;
signal global_clk_c : std_logic;
signal \ctrl_idcodeArea_shifter_25\ : std_logic;
signal \ctrl_idcodeArea_shifter_24\ : std_logic;
signal \ctrl_idcodeArea_shifter_27\ : std_logic;
signal \ctrl_idcodeArea_shifter_26\ : std_logic;
signal io_jtag_tdi_c : std_logic;
signal \ctrl_idcodeArea_shifter_23\ : std_logic;
signal \ctrl_idcodeArea_shifter_22\ : std_logic;
signal \ctrl_idcodeArea_shifter_21\ : std_logic;
signal \ctrl_idcodeArea_shifter_18\ : std_logic;
signal n15 : std_logic;
signal \ctrl_idcodeArea_shifter_20\ : std_logic;
signal n1489 : std_logic;
signal \ctrl_idcodeArea_shifter_19\ : std_logic;
signal \n17_cascade_\ : std_logic;
signal \n1687_cascade_\ : std_logic;
signal n2234 : std_logic;
signal n8 : std_logic;
signal n2198 : std_logic;
signal \ctrl_tap_instructionShift_0\ : std_logic;
signal ctrl_tap_bypass : std_logic;
signal \n2198_cascade_\ : std_logic;
signal n4 : std_logic;
signal \ctrl_tap_tdoUnbufferd_N_213\ : std_logic;
signal n1686 : std_logic;
signal \n112_cascade_\ : std_logic;
signal n929 : std_logic;
signal n1117 : std_logic;
signal \n2260_cascade_\ : std_logic;
signal n1119 : std_logic;
signal ctrl_tap_fsm_state_3 : std_logic;
signal ctrl_tap_fsm_state_2 : std_logic;
signal \ctrl_tap_fsm_stateNext_3__N_10_c_3\ : std_logic;
signal ctrl_tap_fsm_state_1 : std_logic;
signal n2243 : std_logic;
signal n2186 : std_logic;
signal ctrl_tap_fsm_state_0 : std_logic;
signal io_leds_c_1 : std_logic;
signal \ctrl_ledsArea_shifter_1\ : std_logic;
signal \ctrl_ledsArea_store_3\ : std_logic;
signal \ctrl_ledsArea_shifter_3\ : std_logic;
signal io_leds_c_5 : std_logic;
signal \ctrl_ledsArea_shifter_5\ : std_logic;
signal \ctrl_ledsArea_shifter_7\ : std_logic;
signal n1638 : std_logic;
signal io_leds_c_6 : std_logic;
signal n7_adj_2 : std_logic;
signal \ctrl_ledsArea_shifter_6\ : std_logic;
signal n1275 : std_logic;
signal \ctrl_ledsArea_shifter_4\ : std_logic;
signal io_leds_c_4 : std_logic;
signal \ctrl_ledsArea_shifter_2\ : std_logic;
signal n2110 : std_logic;
signal io_leds_c_2 : std_logic;
signal io_jtag_tck_c : std_logic;
signal \_gnd_net_\ : std_logic;

signal global_clk_wire : std_logic;
signal io_jtag_tms_wire : std_logic;
signal global_reset_wire : std_logic;
signal io_jtag_tdi_wire : std_logic;
signal io_jtag_tdo_wire : std_logic;
signal io_leds_wire : std_logic_vector(7 downto 0);
signal io_jtag_tck_wire : std_logic;

begin
    global_clk_wire <= global_clk;
    io_jtag_tms_wire <= io_jtag_tms;
    global_reset_wire <= global_reset;
    io_jtag_tdi_wire <= io_jtag_tdi;
    io_jtag_tdo <= io_jtag_tdo_wire;
    io_leds <= io_leds_wire;
    io_jtag_tck_wire <= io_jtag_tck;

    \global_clk_pad_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__4908\,
            GLOBALBUFFEROUTPUT => global_clk_c
        );

    \global_clk_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4910\,
            DIN => \N__4909\,
            DOUT => \N__4908\,
            PACKAGEPIN => global_clk_wire
        );

    \global_clk_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__4910\,
            PADOUT => \N__4909\,
            PADIN => \N__4908\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \ctrl_tap_fsm_stateNext_3__N_10_pad_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4899\,
            DIN => \N__4898\,
            DOUT => \N__4897\,
            PACKAGEPIN => io_jtag_tms_wire
        );

    \ctrl_tap_fsm_stateNext_3__N_10_pad_3_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__4899\,
            PADOUT => \N__4898\,
            PADIN => \N__4897\,
            CLOCKENABLE => 'H',
            DIN0 => \ctrl_tap_fsm_stateNext_3__N_10_c_3\,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \global_reset_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4890\,
            DIN => \N__4889\,
            DOUT => \N__4888\,
            PACKAGEPIN => global_reset_wire
        );

    \global_reset_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__4890\,
            PADOUT => \N__4889\,
            PADIN => \N__4888\,
            CLOCKENABLE => 'H',
            DIN0 => global_reset_c,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \io_jtag_tdi_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4881\,
            DIN => \N__4880\,
            DOUT => \N__4879\,
            PACKAGEPIN => io_jtag_tdi_wire
        );

    \io_jtag_tdi_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__4881\,
            PADOUT => \N__4880\,
            PADIN => \N__4879\,
            CLOCKENABLE => 'H',
            DIN0 => io_jtag_tdi_c,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \io_jtag_tdo_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4872\,
            DIN => \N__4871\,
            DOUT => \N__4870\,
            PACKAGEPIN => io_jtag_tdo_wire
        );

    \io_jtag_tdo_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "010101",
            NEG_TRIGGER => '1'
        )
    port map (
            PADOEN => \N__4872\,
            PADOUT => \N__4871\,
            PADIN => \N__4870\,
            CLOCKENABLE => \VCCG0\,
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__2246\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => \N__4322\,
            OUTPUTENABLE => '0'
        );

    \io_leds_pad_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4863\,
            DIN => \N__4862\,
            DOUT => \N__4861\,
            PACKAGEPIN => io_leds_wire(0)
        );

    \io_leds_pad_0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__4863\,
            PADOUT => \N__4862\,
            PADIN => \N__4861\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__1892\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \io_leds_pad_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4854\,
            DIN => \N__4853\,
            DOUT => \N__4852\,
            PACKAGEPIN => io_leds_wire(1)
        );

    \io_leds_pad_1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__4854\,
            PADOUT => \N__4853\,
            PADIN => \N__4852\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__4772\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \io_leds_pad_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4845\,
            DIN => \N__4844\,
            DOUT => \N__4843\,
            PACKAGEPIN => io_leds_wire(2)
        );

    \io_leds_pad_2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__4845\,
            PADOUT => \N__4844\,
            PADIN => \N__4843\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__4355\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \io_leds_pad_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4836\,
            DIN => \N__4835\,
            DOUT => \N__4834\,
            PACKAGEPIN => io_leds_wire(3)
        );

    \io_leds_pad_3_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__4836\,
            PADOUT => \N__4835\,
            PADIN => \N__4834\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__2864\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \io_leds_pad_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4827\,
            DIN => \N__4826\,
            DOUT => \N__4825\,
            PACKAGEPIN => io_leds_wire(4)
        );

    \io_leds_pad_4_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__4827\,
            PADOUT => \N__4826\,
            PADIN => \N__4825\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__4457\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \io_leds_pad_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4818\,
            DIN => \N__4817\,
            DOUT => \N__4816\,
            PACKAGEPIN => io_leds_wire(5)
        );

    \io_leds_pad_5_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__4818\,
            PADOUT => \N__4817\,
            PADIN => \N__4816\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__4697\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \io_leds_pad_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4809\,
            DIN => \N__4808\,
            DOUT => \N__4807\,
            PACKAGEPIN => io_leds_wire(6)
        );

    \io_leds_pad_6_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__4809\,
            PADOUT => \N__4808\,
            PADIN => \N__4807\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__4607\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \io_leds_pad_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4800\,
            DIN => \N__4799\,
            DOUT => \N__4798\,
            PACKAGEPIN => io_leds_wire(7)
        );

    \io_leds_pad_7_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__4800\,
            PADOUT => \N__4799\,
            PADIN => \N__4798\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__2807\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \io_jtag_tck_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4791\,
            DIN => \N__4790\,
            DOUT => \N__4789\,
            PACKAGEPIN => io_jtag_tck_wire
        );

    \io_jtag_tck_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__4791\,
            PADOUT => \N__4790\,
            PADIN => \N__4789\,
            CLOCKENABLE => 'H',
            DIN0 => io_jtag_tck_pad_gb_input,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \I__1134\ : IoInMux
    port map (
            O => \N__4772\,
            I => \N__4769\
        );

    \I__1133\ : LocalMux
    port map (
            O => \N__4769\,
            I => \N__4766\
        );

    \I__1132\ : IoSpan4Mux
    port map (
            O => \N__4766\,
            I => \N__4763\
        );

    \I__1131\ : Span4Mux_s2_h
    port map (
            O => \N__4763\,
            I => \N__4759\
        );

    \I__1130\ : CascadeMux
    port map (
            O => \N__4762\,
            I => \N__4756\
        );

    \I__1129\ : Span4Mux_h
    port map (
            O => \N__4759\,
            I => \N__4752\
        );

    \I__1128\ : InMux
    port map (
            O => \N__4756\,
            I => \N__4749\
        );

    \I__1127\ : InMux
    port map (
            O => \N__4755\,
            I => \N__4746\
        );

    \I__1126\ : Odrv4
    port map (
            O => \N__4752\,
            I => io_leds_c_1
        );

    \I__1125\ : LocalMux
    port map (
            O => \N__4749\,
            I => io_leds_c_1
        );

    \I__1124\ : LocalMux
    port map (
            O => \N__4746\,
            I => io_leds_c_1
        );

    \I__1123\ : InMux
    port map (
            O => \N__4739\,
            I => \N__4735\
        );

    \I__1122\ : InMux
    port map (
            O => \N__4738\,
            I => \N__4732\
        );

    \I__1121\ : LocalMux
    port map (
            O => \N__4735\,
            I => \N__4729\
        );

    \I__1120\ : LocalMux
    port map (
            O => \N__4732\,
            I => \ctrl_ledsArea_shifter_1\
        );

    \I__1119\ : Odrv12
    port map (
            O => \N__4729\,
            I => \ctrl_ledsArea_shifter_1\
        );

    \I__1118\ : CascadeMux
    port map (
            O => \N__4724\,
            I => \N__4721\
        );

    \I__1117\ : InMux
    port map (
            O => \N__4721\,
            I => \N__4717\
        );

    \I__1116\ : InMux
    port map (
            O => \N__4720\,
            I => \N__4714\
        );

    \I__1115\ : LocalMux
    port map (
            O => \N__4717\,
            I => \ctrl_ledsArea_store_3\
        );

    \I__1114\ : LocalMux
    port map (
            O => \N__4714\,
            I => \ctrl_ledsArea_store_3\
        );

    \I__1113\ : InMux
    port map (
            O => \N__4709\,
            I => \N__4705\
        );

    \I__1112\ : InMux
    port map (
            O => \N__4708\,
            I => \N__4702\
        );

    \I__1111\ : LocalMux
    port map (
            O => \N__4705\,
            I => \ctrl_ledsArea_shifter_3\
        );

    \I__1110\ : LocalMux
    port map (
            O => \N__4702\,
            I => \ctrl_ledsArea_shifter_3\
        );

    \I__1109\ : IoInMux
    port map (
            O => \N__4697\,
            I => \N__4693\
        );

    \I__1108\ : CascadeMux
    port map (
            O => \N__4696\,
            I => \N__4690\
        );

    \I__1107\ : LocalMux
    port map (
            O => \N__4693\,
            I => \N__4687\
        );

    \I__1106\ : InMux
    port map (
            O => \N__4690\,
            I => \N__4684\
        );

    \I__1105\ : IoSpan4Mux
    port map (
            O => \N__4687\,
            I => \N__4681\
        );

    \I__1104\ : LocalMux
    port map (
            O => \N__4684\,
            I => \N__4678\
        );

    \I__1103\ : Span4Mux_s3_h
    port map (
            O => \N__4681\,
            I => \N__4672\
        );

    \I__1102\ : Span4Mux_v
    port map (
            O => \N__4678\,
            I => \N__4672\
        );

    \I__1101\ : InMux
    port map (
            O => \N__4677\,
            I => \N__4669\
        );

    \I__1100\ : Odrv4
    port map (
            O => \N__4672\,
            I => io_leds_c_5
        );

    \I__1099\ : LocalMux
    port map (
            O => \N__4669\,
            I => io_leds_c_5
        );

    \I__1098\ : InMux
    port map (
            O => \N__4664\,
            I => \N__4660\
        );

    \I__1097\ : CascadeMux
    port map (
            O => \N__4663\,
            I => \N__4657\
        );

    \I__1096\ : LocalMux
    port map (
            O => \N__4660\,
            I => \N__4654\
        );

    \I__1095\ : InMux
    port map (
            O => \N__4657\,
            I => \N__4651\
        );

    \I__1094\ : Span4Mux_h
    port map (
            O => \N__4654\,
            I => \N__4648\
        );

    \I__1093\ : LocalMux
    port map (
            O => \N__4651\,
            I => \ctrl_ledsArea_shifter_5\
        );

    \I__1092\ : Odrv4
    port map (
            O => \N__4648\,
            I => \ctrl_ledsArea_shifter_5\
        );

    \I__1091\ : InMux
    port map (
            O => \N__4643\,
            I => \N__4639\
        );

    \I__1090\ : InMux
    port map (
            O => \N__4642\,
            I => \N__4636\
        );

    \I__1089\ : LocalMux
    port map (
            O => \N__4639\,
            I => \N__4633\
        );

    \I__1088\ : LocalMux
    port map (
            O => \N__4636\,
            I => \ctrl_ledsArea_shifter_7\
        );

    \I__1087\ : Odrv12
    port map (
            O => \N__4633\,
            I => \ctrl_ledsArea_shifter_7\
        );

    \I__1086\ : InMux
    port map (
            O => \N__4628\,
            I => \N__4619\
        );

    \I__1085\ : InMux
    port map (
            O => \N__4627\,
            I => \N__4619\
        );

    \I__1084\ : InMux
    port map (
            O => \N__4626\,
            I => \N__4612\
        );

    \I__1083\ : InMux
    port map (
            O => \N__4625\,
            I => \N__4612\
        );

    \I__1082\ : InMux
    port map (
            O => \N__4624\,
            I => \N__4612\
        );

    \I__1081\ : LocalMux
    port map (
            O => \N__4619\,
            I => n1638
        );

    \I__1080\ : LocalMux
    port map (
            O => \N__4612\,
            I => n1638
        );

    \I__1079\ : IoInMux
    port map (
            O => \N__4607\,
            I => \N__4604\
        );

    \I__1078\ : LocalMux
    port map (
            O => \N__4604\,
            I => \N__4601\
        );

    \I__1077\ : IoSpan4Mux
    port map (
            O => \N__4601\,
            I => \N__4597\
        );

    \I__1076\ : CascadeMux
    port map (
            O => \N__4600\,
            I => \N__4594\
        );

    \I__1075\ : Span4Mux_s0_h
    port map (
            O => \N__4597\,
            I => \N__4591\
        );

    \I__1074\ : InMux
    port map (
            O => \N__4594\,
            I => \N__4588\
        );

    \I__1073\ : Span4Mux_h
    port map (
            O => \N__4591\,
            I => \N__4583\
        );

    \I__1072\ : LocalMux
    port map (
            O => \N__4588\,
            I => \N__4583\
        );

    \I__1071\ : Span4Mux_h
    port map (
            O => \N__4583\,
            I => \N__4579\
        );

    \I__1070\ : InMux
    port map (
            O => \N__4582\,
            I => \N__4576\
        );

    \I__1069\ : Odrv4
    port map (
            O => \N__4579\,
            I => io_leds_c_6
        );

    \I__1068\ : LocalMux
    port map (
            O => \N__4576\,
            I => io_leds_c_6
        );

    \I__1067\ : InMux
    port map (
            O => \N__4571\,
            I => \N__4567\
        );

    \I__1066\ : InMux
    port map (
            O => \N__4570\,
            I => \N__4564\
        );

    \I__1065\ : LocalMux
    port map (
            O => \N__4567\,
            I => \N__4561\
        );

    \I__1064\ : LocalMux
    port map (
            O => \N__4564\,
            I => \N__4558\
        );

    \I__1063\ : Span4Mux_v
    port map (
            O => \N__4561\,
            I => \N__4548\
        );

    \I__1062\ : Span4Mux_v
    port map (
            O => \N__4558\,
            I => \N__4545\
        );

    \I__1061\ : InMux
    port map (
            O => \N__4557\,
            I => \N__4534\
        );

    \I__1060\ : InMux
    port map (
            O => \N__4556\,
            I => \N__4534\
        );

    \I__1059\ : InMux
    port map (
            O => \N__4555\,
            I => \N__4534\
        );

    \I__1058\ : InMux
    port map (
            O => \N__4554\,
            I => \N__4534\
        );

    \I__1057\ : InMux
    port map (
            O => \N__4553\,
            I => \N__4534\
        );

    \I__1056\ : InMux
    port map (
            O => \N__4552\,
            I => \N__4529\
        );

    \I__1055\ : InMux
    port map (
            O => \N__4551\,
            I => \N__4529\
        );

    \I__1054\ : Odrv4
    port map (
            O => \N__4548\,
            I => n7_adj_2
        );

    \I__1053\ : Odrv4
    port map (
            O => \N__4545\,
            I => n7_adj_2
        );

    \I__1052\ : LocalMux
    port map (
            O => \N__4534\,
            I => n7_adj_2
        );

    \I__1051\ : LocalMux
    port map (
            O => \N__4529\,
            I => n7_adj_2
        );

    \I__1050\ : InMux
    port map (
            O => \N__4520\,
            I => \N__4517\
        );

    \I__1049\ : LocalMux
    port map (
            O => \N__4517\,
            I => \N__4514\
        );

    \I__1048\ : Span4Mux_h
    port map (
            O => \N__4514\,
            I => \N__4510\
        );

    \I__1047\ : InMux
    port map (
            O => \N__4513\,
            I => \N__4507\
        );

    \I__1046\ : Odrv4
    port map (
            O => \N__4510\,
            I => \ctrl_ledsArea_shifter_6\
        );

    \I__1045\ : LocalMux
    port map (
            O => \N__4507\,
            I => \ctrl_ledsArea_shifter_6\
        );

    \I__1044\ : CEMux
    port map (
            O => \N__4502\,
            I => \N__4499\
        );

    \I__1043\ : LocalMux
    port map (
            O => \N__4499\,
            I => \N__4494\
        );

    \I__1042\ : CEMux
    port map (
            O => \N__4498\,
            I => \N__4491\
        );

    \I__1041\ : CEMux
    port map (
            O => \N__4497\,
            I => \N__4488\
        );

    \I__1040\ : Span4Mux_h
    port map (
            O => \N__4494\,
            I => \N__4485\
        );

    \I__1039\ : LocalMux
    port map (
            O => \N__4491\,
            I => \N__4482\
        );

    \I__1038\ : LocalMux
    port map (
            O => \N__4488\,
            I => \N__4479\
        );

    \I__1037\ : Odrv4
    port map (
            O => \N__4485\,
            I => n1275
        );

    \I__1036\ : Odrv4
    port map (
            O => \N__4482\,
            I => n1275
        );

    \I__1035\ : Odrv4
    port map (
            O => \N__4479\,
            I => n1275
        );

    \I__1034\ : InMux
    port map (
            O => \N__4472\,
            I => \N__4468\
        );

    \I__1033\ : InMux
    port map (
            O => \N__4471\,
            I => \N__4465\
        );

    \I__1032\ : LocalMux
    port map (
            O => \N__4468\,
            I => \N__4462\
        );

    \I__1031\ : LocalMux
    port map (
            O => \N__4465\,
            I => \ctrl_ledsArea_shifter_4\
        );

    \I__1030\ : Odrv4
    port map (
            O => \N__4462\,
            I => \ctrl_ledsArea_shifter_4\
        );

    \I__1029\ : IoInMux
    port map (
            O => \N__4457\,
            I => \N__4454\
        );

    \I__1028\ : LocalMux
    port map (
            O => \N__4454\,
            I => \N__4451\
        );

    \I__1027\ : Span12Mux_s5_h
    port map (
            O => \N__4451\,
            I => \N__4446\
        );

    \I__1026\ : InMux
    port map (
            O => \N__4450\,
            I => \N__4443\
        );

    \I__1025\ : InMux
    port map (
            O => \N__4449\,
            I => \N__4440\
        );

    \I__1024\ : Odrv12
    port map (
            O => \N__4446\,
            I => io_leds_c_4
        );

    \I__1023\ : LocalMux
    port map (
            O => \N__4443\,
            I => io_leds_c_4
        );

    \I__1022\ : LocalMux
    port map (
            O => \N__4440\,
            I => io_leds_c_4
        );

    \I__1021\ : InMux
    port map (
            O => \N__4433\,
            I => \N__4430\
        );

    \I__1020\ : LocalMux
    port map (
            O => \N__4430\,
            I => \N__4426\
        );

    \I__1019\ : InMux
    port map (
            O => \N__4429\,
            I => \N__4423\
        );

    \I__1018\ : Odrv4
    port map (
            O => \N__4426\,
            I => \ctrl_ledsArea_shifter_2\
        );

    \I__1017\ : LocalMux
    port map (
            O => \N__4423\,
            I => \ctrl_ledsArea_shifter_2\
        );

    \I__1016\ : InMux
    port map (
            O => \N__4418\,
            I => \N__4411\
        );

    \I__1015\ : InMux
    port map (
            O => \N__4417\,
            I => \N__4408\
        );

    \I__1014\ : InMux
    port map (
            O => \N__4416\,
            I => \N__4405\
        );

    \I__1013\ : InMux
    port map (
            O => \N__4415\,
            I => \N__4402\
        );

    \I__1012\ : InMux
    port map (
            O => \N__4414\,
            I => \N__4397\
        );

    \I__1011\ : LocalMux
    port map (
            O => \N__4411\,
            I => \N__4394\
        );

    \I__1010\ : LocalMux
    port map (
            O => \N__4408\,
            I => \N__4388\
        );

    \I__1009\ : LocalMux
    port map (
            O => \N__4405\,
            I => \N__4388\
        );

    \I__1008\ : LocalMux
    port map (
            O => \N__4402\,
            I => \N__4385\
        );

    \I__1007\ : InMux
    port map (
            O => \N__4401\,
            I => \N__4380\
        );

    \I__1006\ : InMux
    port map (
            O => \N__4400\,
            I => \N__4380\
        );

    \I__1005\ : LocalMux
    port map (
            O => \N__4397\,
            I => \N__4377\
        );

    \I__1004\ : Span4Mux_h
    port map (
            O => \N__4394\,
            I => \N__4374\
        );

    \I__1003\ : InMux
    port map (
            O => \N__4393\,
            I => \N__4371\
        );

    \I__1002\ : Span4Mux_v
    port map (
            O => \N__4388\,
            I => \N__4364\
        );

    \I__1001\ : Span4Mux_v
    port map (
            O => \N__4385\,
            I => \N__4364\
        );

    \I__1000\ : LocalMux
    port map (
            O => \N__4380\,
            I => \N__4364\
        );

    \I__999\ : Odrv4
    port map (
            O => \N__4377\,
            I => n2110
        );

    \I__998\ : Odrv4
    port map (
            O => \N__4374\,
            I => n2110
        );

    \I__997\ : LocalMux
    port map (
            O => \N__4371\,
            I => n2110
        );

    \I__996\ : Odrv4
    port map (
            O => \N__4364\,
            I => n2110
        );

    \I__995\ : IoInMux
    port map (
            O => \N__4355\,
            I => \N__4352\
        );

    \I__994\ : LocalMux
    port map (
            O => \N__4352\,
            I => \N__4348\
        );

    \I__993\ : CascadeMux
    port map (
            O => \N__4351\,
            I => \N__4345\
        );

    \I__992\ : IoSpan4Mux
    port map (
            O => \N__4348\,
            I => \N__4342\
        );

    \I__991\ : InMux
    port map (
            O => \N__4345\,
            I => \N__4339\
        );

    \I__990\ : Span4Mux_s2_h
    port map (
            O => \N__4342\,
            I => \N__4335\
        );

    \I__989\ : LocalMux
    port map (
            O => \N__4339\,
            I => \N__4332\
        );

    \I__988\ : InMux
    port map (
            O => \N__4338\,
            I => \N__4329\
        );

    \I__987\ : Odrv4
    port map (
            O => \N__4335\,
            I => io_leds_c_2
        );

    \I__986\ : Odrv4
    port map (
            O => \N__4332\,
            I => io_leds_c_2
        );

    \I__985\ : LocalMux
    port map (
            O => \N__4329\,
            I => io_leds_c_2
        );

    \I__984\ : ClkMux
    port map (
            O => \N__4322\,
            I => \N__4265\
        );

    \I__983\ : ClkMux
    port map (
            O => \N__4321\,
            I => \N__4265\
        );

    \I__982\ : ClkMux
    port map (
            O => \N__4320\,
            I => \N__4265\
        );

    \I__981\ : ClkMux
    port map (
            O => \N__4319\,
            I => \N__4265\
        );

    \I__980\ : ClkMux
    port map (
            O => \N__4318\,
            I => \N__4265\
        );

    \I__979\ : ClkMux
    port map (
            O => \N__4317\,
            I => \N__4265\
        );

    \I__978\ : ClkMux
    port map (
            O => \N__4316\,
            I => \N__4265\
        );

    \I__977\ : ClkMux
    port map (
            O => \N__4315\,
            I => \N__4265\
        );

    \I__976\ : ClkMux
    port map (
            O => \N__4314\,
            I => \N__4265\
        );

    \I__975\ : ClkMux
    port map (
            O => \N__4313\,
            I => \N__4265\
        );

    \I__974\ : ClkMux
    port map (
            O => \N__4312\,
            I => \N__4265\
        );

    \I__973\ : ClkMux
    port map (
            O => \N__4311\,
            I => \N__4265\
        );

    \I__972\ : ClkMux
    port map (
            O => \N__4310\,
            I => \N__4265\
        );

    \I__971\ : ClkMux
    port map (
            O => \N__4309\,
            I => \N__4265\
        );

    \I__970\ : ClkMux
    port map (
            O => \N__4308\,
            I => \N__4265\
        );

    \I__969\ : ClkMux
    port map (
            O => \N__4307\,
            I => \N__4265\
        );

    \I__968\ : ClkMux
    port map (
            O => \N__4306\,
            I => \N__4265\
        );

    \I__967\ : ClkMux
    port map (
            O => \N__4305\,
            I => \N__4265\
        );

    \I__966\ : ClkMux
    port map (
            O => \N__4304\,
            I => \N__4265\
        );

    \I__965\ : GlobalMux
    port map (
            O => \N__4265\,
            I => \N__4262\
        );

    \I__964\ : gio2CtrlBuf
    port map (
            O => \N__4262\,
            I => io_jtag_tck_c
        );

    \I__963\ : InMux
    port map (
            O => \N__4259\,
            I => \N__4255\
        );

    \I__962\ : InMux
    port map (
            O => \N__4258\,
            I => \N__4252\
        );

    \I__961\ : LocalMux
    port map (
            O => \N__4255\,
            I => n1686
        );

    \I__960\ : LocalMux
    port map (
            O => \N__4252\,
            I => n1686
        );

    \I__959\ : CascadeMux
    port map (
            O => \N__4247\,
            I => \n112_cascade_\
        );

    \I__958\ : InMux
    port map (
            O => \N__4244\,
            I => \N__4241\
        );

    \I__957\ : LocalMux
    port map (
            O => \N__4241\,
            I => \N__4238\
        );

    \I__956\ : Odrv4
    port map (
            O => \N__4238\,
            I => n929
        );

    \I__955\ : CascadeMux
    port map (
            O => \N__4235\,
            I => \N__4232\
        );

    \I__954\ : InMux
    port map (
            O => \N__4232\,
            I => \N__4228\
        );

    \I__953\ : InMux
    port map (
            O => \N__4231\,
            I => \N__4223\
        );

    \I__952\ : LocalMux
    port map (
            O => \N__4228\,
            I => \N__4220\
        );

    \I__951\ : InMux
    port map (
            O => \N__4227\,
            I => \N__4215\
        );

    \I__950\ : InMux
    port map (
            O => \N__4226\,
            I => \N__4215\
        );

    \I__949\ : LocalMux
    port map (
            O => \N__4223\,
            I => n1117
        );

    \I__948\ : Odrv4
    port map (
            O => \N__4220\,
            I => n1117
        );

    \I__947\ : LocalMux
    port map (
            O => \N__4215\,
            I => n1117
        );

    \I__946\ : CascadeMux
    port map (
            O => \N__4208\,
            I => \n2260_cascade_\
        );

    \I__945\ : InMux
    port map (
            O => \N__4205\,
            I => \N__4195\
        );

    \I__944\ : InMux
    port map (
            O => \N__4204\,
            I => \N__4192\
        );

    \I__943\ : InMux
    port map (
            O => \N__4203\,
            I => \N__4189\
        );

    \I__942\ : InMux
    port map (
            O => \N__4202\,
            I => \N__4184\
        );

    \I__941\ : InMux
    port map (
            O => \N__4201\,
            I => \N__4184\
        );

    \I__940\ : InMux
    port map (
            O => \N__4200\,
            I => \N__4181\
        );

    \I__939\ : InMux
    port map (
            O => \N__4199\,
            I => \N__4178\
        );

    \I__938\ : InMux
    port map (
            O => \N__4198\,
            I => \N__4175\
        );

    \I__937\ : LocalMux
    port map (
            O => \N__4195\,
            I => n1119
        );

    \I__936\ : LocalMux
    port map (
            O => \N__4192\,
            I => n1119
        );

    \I__935\ : LocalMux
    port map (
            O => \N__4189\,
            I => n1119
        );

    \I__934\ : LocalMux
    port map (
            O => \N__4184\,
            I => n1119
        );

    \I__933\ : LocalMux
    port map (
            O => \N__4181\,
            I => n1119
        );

    \I__932\ : LocalMux
    port map (
            O => \N__4178\,
            I => n1119
        );

    \I__931\ : LocalMux
    port map (
            O => \N__4175\,
            I => n1119
        );

    \I__930\ : CascadeMux
    port map (
            O => \N__4160\,
            I => \N__4157\
        );

    \I__929\ : InMux
    port map (
            O => \N__4157\,
            I => \N__4145\
        );

    \I__928\ : InMux
    port map (
            O => \N__4156\,
            I => \N__4145\
        );

    \I__927\ : InMux
    port map (
            O => \N__4155\,
            I => \N__4145\
        );

    \I__926\ : CascadeMux
    port map (
            O => \N__4154\,
            I => \N__4137\
        );

    \I__925\ : InMux
    port map (
            O => \N__4153\,
            I => \N__4134\
        );

    \I__924\ : InMux
    port map (
            O => \N__4152\,
            I => \N__4131\
        );

    \I__923\ : LocalMux
    port map (
            O => \N__4145\,
            I => \N__4128\
        );

    \I__922\ : CascadeMux
    port map (
            O => \N__4144\,
            I => \N__4125\
        );

    \I__921\ : CascadeMux
    port map (
            O => \N__4143\,
            I => \N__4117\
        );

    \I__920\ : InMux
    port map (
            O => \N__4142\,
            I => \N__4107\
        );

    \I__919\ : InMux
    port map (
            O => \N__4141\,
            I => \N__4100\
        );

    \I__918\ : InMux
    port map (
            O => \N__4140\,
            I => \N__4100\
        );

    \I__917\ : InMux
    port map (
            O => \N__4137\,
            I => \N__4100\
        );

    \I__916\ : LocalMux
    port map (
            O => \N__4134\,
            I => \N__4095\
        );

    \I__915\ : LocalMux
    port map (
            O => \N__4131\,
            I => \N__4095\
        );

    \I__914\ : Span4Mux_v
    port map (
            O => \N__4128\,
            I => \N__4092\
        );

    \I__913\ : InMux
    port map (
            O => \N__4125\,
            I => \N__4083\
        );

    \I__912\ : InMux
    port map (
            O => \N__4124\,
            I => \N__4083\
        );

    \I__911\ : InMux
    port map (
            O => \N__4123\,
            I => \N__4083\
        );

    \I__910\ : InMux
    port map (
            O => \N__4122\,
            I => \N__4083\
        );

    \I__909\ : InMux
    port map (
            O => \N__4121\,
            I => \N__4076\
        );

    \I__908\ : InMux
    port map (
            O => \N__4120\,
            I => \N__4076\
        );

    \I__907\ : InMux
    port map (
            O => \N__4117\,
            I => \N__4076\
        );

    \I__906\ : InMux
    port map (
            O => \N__4116\,
            I => \N__4067\
        );

    \I__905\ : InMux
    port map (
            O => \N__4115\,
            I => \N__4067\
        );

    \I__904\ : InMux
    port map (
            O => \N__4114\,
            I => \N__4067\
        );

    \I__903\ : InMux
    port map (
            O => \N__4113\,
            I => \N__4067\
        );

    \I__902\ : InMux
    port map (
            O => \N__4112\,
            I => \N__4060\
        );

    \I__901\ : InMux
    port map (
            O => \N__4111\,
            I => \N__4060\
        );

    \I__900\ : InMux
    port map (
            O => \N__4110\,
            I => \N__4060\
        );

    \I__899\ : LocalMux
    port map (
            O => \N__4107\,
            I => ctrl_tap_fsm_state_3
        );

    \I__898\ : LocalMux
    port map (
            O => \N__4100\,
            I => ctrl_tap_fsm_state_3
        );

    \I__897\ : Odrv4
    port map (
            O => \N__4095\,
            I => ctrl_tap_fsm_state_3
        );

    \I__896\ : Odrv4
    port map (
            O => \N__4092\,
            I => ctrl_tap_fsm_state_3
        );

    \I__895\ : LocalMux
    port map (
            O => \N__4083\,
            I => ctrl_tap_fsm_state_3
        );

    \I__894\ : LocalMux
    port map (
            O => \N__4076\,
            I => ctrl_tap_fsm_state_3
        );

    \I__893\ : LocalMux
    port map (
            O => \N__4067\,
            I => ctrl_tap_fsm_state_3
        );

    \I__892\ : LocalMux
    port map (
            O => \N__4060\,
            I => ctrl_tap_fsm_state_3
        );

    \I__891\ : CascadeMux
    port map (
            O => \N__4043\,
            I => \N__4029\
        );

    \I__890\ : CascadeMux
    port map (
            O => \N__4042\,
            I => \N__4024\
        );

    \I__889\ : CascadeMux
    port map (
            O => \N__4041\,
            I => \N__4018\
        );

    \I__888\ : InMux
    port map (
            O => \N__4040\,
            I => \N__4010\
        );

    \I__887\ : InMux
    port map (
            O => \N__4039\,
            I => \N__4010\
        );

    \I__886\ : InMux
    port map (
            O => \N__4038\,
            I => \N__4010\
        );

    \I__885\ : InMux
    port map (
            O => \N__4037\,
            I => \N__4007\
        );

    \I__884\ : InMux
    port map (
            O => \N__4036\,
            I => \N__4004\
        );

    \I__883\ : InMux
    port map (
            O => \N__4035\,
            I => \N__4001\
        );

    \I__882\ : InMux
    port map (
            O => \N__4034\,
            I => \N__3996\
        );

    \I__881\ : InMux
    port map (
            O => \N__4033\,
            I => \N__3996\
        );

    \I__880\ : InMux
    port map (
            O => \N__4032\,
            I => \N__3987\
        );

    \I__879\ : InMux
    port map (
            O => \N__4029\,
            I => \N__3987\
        );

    \I__878\ : InMux
    port map (
            O => \N__4028\,
            I => \N__3987\
        );

    \I__877\ : InMux
    port map (
            O => \N__4027\,
            I => \N__3987\
        );

    \I__876\ : InMux
    port map (
            O => \N__4024\,
            I => \N__3980\
        );

    \I__875\ : InMux
    port map (
            O => \N__4023\,
            I => \N__3980\
        );

    \I__874\ : InMux
    port map (
            O => \N__4022\,
            I => \N__3980\
        );

    \I__873\ : InMux
    port map (
            O => \N__4021\,
            I => \N__3973\
        );

    \I__872\ : InMux
    port map (
            O => \N__4018\,
            I => \N__3973\
        );

    \I__871\ : InMux
    port map (
            O => \N__4017\,
            I => \N__3973\
        );

    \I__870\ : LocalMux
    port map (
            O => \N__4010\,
            I => ctrl_tap_fsm_state_2
        );

    \I__869\ : LocalMux
    port map (
            O => \N__4007\,
            I => ctrl_tap_fsm_state_2
        );

    \I__868\ : LocalMux
    port map (
            O => \N__4004\,
            I => ctrl_tap_fsm_state_2
        );

    \I__867\ : LocalMux
    port map (
            O => \N__4001\,
            I => ctrl_tap_fsm_state_2
        );

    \I__866\ : LocalMux
    port map (
            O => \N__3996\,
            I => ctrl_tap_fsm_state_2
        );

    \I__865\ : LocalMux
    port map (
            O => \N__3987\,
            I => ctrl_tap_fsm_state_2
        );

    \I__864\ : LocalMux
    port map (
            O => \N__3980\,
            I => ctrl_tap_fsm_state_2
        );

    \I__863\ : LocalMux
    port map (
            O => \N__3973\,
            I => ctrl_tap_fsm_state_2
        );

    \I__862\ : CascadeMux
    port map (
            O => \N__3956\,
            I => \N__3946\
        );

    \I__861\ : CascadeMux
    port map (
            O => \N__3955\,
            I => \N__3940\
        );

    \I__860\ : InMux
    port map (
            O => \N__3954\,
            I => \N__3934\
        );

    \I__859\ : InMux
    port map (
            O => \N__3953\,
            I => \N__3934\
        );

    \I__858\ : InMux
    port map (
            O => \N__3952\,
            I => \N__3931\
        );

    \I__857\ : InMux
    port map (
            O => \N__3951\,
            I => \N__3926\
        );

    \I__856\ : InMux
    port map (
            O => \N__3950\,
            I => \N__3926\
        );

    \I__855\ : CascadeMux
    port map (
            O => \N__3949\,
            I => \N__3923\
        );

    \I__854\ : InMux
    port map (
            O => \N__3946\,
            I => \N__3920\
        );

    \I__853\ : InMux
    port map (
            O => \N__3945\,
            I => \N__3913\
        );

    \I__852\ : InMux
    port map (
            O => \N__3944\,
            I => \N__3913\
        );

    \I__851\ : InMux
    port map (
            O => \N__3943\,
            I => \N__3913\
        );

    \I__850\ : InMux
    port map (
            O => \N__3940\,
            I => \N__3907\
        );

    \I__849\ : InMux
    port map (
            O => \N__3939\,
            I => \N__3907\
        );

    \I__848\ : LocalMux
    port map (
            O => \N__3934\,
            I => \N__3900\
        );

    \I__847\ : LocalMux
    port map (
            O => \N__3931\,
            I => \N__3900\
        );

    \I__846\ : LocalMux
    port map (
            O => \N__3926\,
            I => \N__3900\
        );

    \I__845\ : InMux
    port map (
            O => \N__3923\,
            I => \N__3897\
        );

    \I__844\ : LocalMux
    port map (
            O => \N__3920\,
            I => \N__3892\
        );

    \I__843\ : LocalMux
    port map (
            O => \N__3913\,
            I => \N__3892\
        );

    \I__842\ : InMux
    port map (
            O => \N__3912\,
            I => \N__3889\
        );

    \I__841\ : LocalMux
    port map (
            O => \N__3907\,
            I => \N__3886\
        );

    \I__840\ : Span4Mux_h
    port map (
            O => \N__3900\,
            I => \N__3883\
        );

    \I__839\ : LocalMux
    port map (
            O => \N__3897\,
            I => \N__3880\
        );

    \I__838\ : Span4Mux_h
    port map (
            O => \N__3892\,
            I => \N__3877\
        );

    \I__837\ : LocalMux
    port map (
            O => \N__3889\,
            I => \N__3874\
        );

    \I__836\ : Span12Mux_s8_h
    port map (
            O => \N__3886\,
            I => \N__3871\
        );

    \I__835\ : Span4Mux_v
    port map (
            O => \N__3883\,
            I => \N__3868\
        );

    \I__834\ : Span4Mux_h
    port map (
            O => \N__3880\,
            I => \N__3865\
        );

    \I__833\ : Span4Mux_v
    port map (
            O => \N__3877\,
            I => \N__3860\
        );

    \I__832\ : Span4Mux_v
    port map (
            O => \N__3874\,
            I => \N__3860\
        );

    \I__831\ : Odrv12
    port map (
            O => \N__3871\,
            I => \ctrl_tap_fsm_stateNext_3__N_10_c_3\
        );

    \I__830\ : Odrv4
    port map (
            O => \N__3868\,
            I => \ctrl_tap_fsm_stateNext_3__N_10_c_3\
        );

    \I__829\ : Odrv4
    port map (
            O => \N__3865\,
            I => \ctrl_tap_fsm_stateNext_3__N_10_c_3\
        );

    \I__828\ : Odrv4
    port map (
            O => \N__3860\,
            I => \ctrl_tap_fsm_stateNext_3__N_10_c_3\
        );

    \I__827\ : CascadeMux
    port map (
            O => \N__3851\,
            I => \N__3844\
        );

    \I__826\ : InMux
    port map (
            O => \N__3850\,
            I => \N__3829\
        );

    \I__825\ : InMux
    port map (
            O => \N__3849\,
            I => \N__3829\
        );

    \I__824\ : InMux
    port map (
            O => \N__3848\,
            I => \N__3829\
        );

    \I__823\ : InMux
    port map (
            O => \N__3847\,
            I => \N__3826\
        );

    \I__822\ : InMux
    port map (
            O => \N__3844\,
            I => \N__3823\
        );

    \I__821\ : InMux
    port map (
            O => \N__3843\,
            I => \N__3807\
        );

    \I__820\ : InMux
    port map (
            O => \N__3842\,
            I => \N__3807\
        );

    \I__819\ : InMux
    port map (
            O => \N__3841\,
            I => \N__3807\
        );

    \I__818\ : InMux
    port map (
            O => \N__3840\,
            I => \N__3804\
        );

    \I__817\ : InMux
    port map (
            O => \N__3839\,
            I => \N__3799\
        );

    \I__816\ : InMux
    port map (
            O => \N__3838\,
            I => \N__3799\
        );

    \I__815\ : InMux
    port map (
            O => \N__3837\,
            I => \N__3794\
        );

    \I__814\ : InMux
    port map (
            O => \N__3836\,
            I => \N__3794\
        );

    \I__813\ : LocalMux
    port map (
            O => \N__3829\,
            I => \N__3791\
        );

    \I__812\ : LocalMux
    port map (
            O => \N__3826\,
            I => \N__3786\
        );

    \I__811\ : LocalMux
    port map (
            O => \N__3823\,
            I => \N__3786\
        );

    \I__810\ : InMux
    port map (
            O => \N__3822\,
            I => \N__3779\
        );

    \I__809\ : InMux
    port map (
            O => \N__3821\,
            I => \N__3779\
        );

    \I__808\ : InMux
    port map (
            O => \N__3820\,
            I => \N__3779\
        );

    \I__807\ : InMux
    port map (
            O => \N__3819\,
            I => \N__3774\
        );

    \I__806\ : InMux
    port map (
            O => \N__3818\,
            I => \N__3774\
        );

    \I__805\ : InMux
    port map (
            O => \N__3817\,
            I => \N__3765\
        );

    \I__804\ : InMux
    port map (
            O => \N__3816\,
            I => \N__3765\
        );

    \I__803\ : InMux
    port map (
            O => \N__3815\,
            I => \N__3765\
        );

    \I__802\ : InMux
    port map (
            O => \N__3814\,
            I => \N__3765\
        );

    \I__801\ : LocalMux
    port map (
            O => \N__3807\,
            I => ctrl_tap_fsm_state_1
        );

    \I__800\ : LocalMux
    port map (
            O => \N__3804\,
            I => ctrl_tap_fsm_state_1
        );

    \I__799\ : LocalMux
    port map (
            O => \N__3799\,
            I => ctrl_tap_fsm_state_1
        );

    \I__798\ : LocalMux
    port map (
            O => \N__3794\,
            I => ctrl_tap_fsm_state_1
        );

    \I__797\ : Odrv4
    port map (
            O => \N__3791\,
            I => ctrl_tap_fsm_state_1
        );

    \I__796\ : Odrv4
    port map (
            O => \N__3786\,
            I => ctrl_tap_fsm_state_1
        );

    \I__795\ : LocalMux
    port map (
            O => \N__3779\,
            I => ctrl_tap_fsm_state_1
        );

    \I__794\ : LocalMux
    port map (
            O => \N__3774\,
            I => ctrl_tap_fsm_state_1
        );

    \I__793\ : LocalMux
    port map (
            O => \N__3765\,
            I => ctrl_tap_fsm_state_1
        );

    \I__792\ : InMux
    port map (
            O => \N__3746\,
            I => \N__3743\
        );

    \I__791\ : LocalMux
    port map (
            O => \N__3743\,
            I => n2243
        );

    \I__790\ : InMux
    port map (
            O => \N__3740\,
            I => \N__3737\
        );

    \I__789\ : LocalMux
    port map (
            O => \N__3737\,
            I => n2186
        );

    \I__788\ : InMux
    port map (
            O => \N__3734\,
            I => \N__3727\
        );

    \I__787\ : CascadeMux
    port map (
            O => \N__3733\,
            I => \N__3716\
        );

    \I__786\ : CascadeMux
    port map (
            O => \N__3732\,
            I => \N__3712\
        );

    \I__785\ : InMux
    port map (
            O => \N__3731\,
            I => \N__3708\
        );

    \I__784\ : CascadeMux
    port map (
            O => \N__3730\,
            I => \N__3700\
        );

    \I__783\ : LocalMux
    port map (
            O => \N__3727\,
            I => \N__3694\
        );

    \I__782\ : InMux
    port map (
            O => \N__3726\,
            I => \N__3689\
        );

    \I__781\ : InMux
    port map (
            O => \N__3725\,
            I => \N__3689\
        );

    \I__780\ : InMux
    port map (
            O => \N__3724\,
            I => \N__3680\
        );

    \I__779\ : InMux
    port map (
            O => \N__3723\,
            I => \N__3680\
        );

    \I__778\ : InMux
    port map (
            O => \N__3722\,
            I => \N__3680\
        );

    \I__777\ : InMux
    port map (
            O => \N__3721\,
            I => \N__3680\
        );

    \I__776\ : InMux
    port map (
            O => \N__3720\,
            I => \N__3677\
        );

    \I__775\ : InMux
    port map (
            O => \N__3719\,
            I => \N__3672\
        );

    \I__774\ : InMux
    port map (
            O => \N__3716\,
            I => \N__3672\
        );

    \I__773\ : InMux
    port map (
            O => \N__3715\,
            I => \N__3669\
        );

    \I__772\ : InMux
    port map (
            O => \N__3712\,
            I => \N__3664\
        );

    \I__771\ : InMux
    port map (
            O => \N__3711\,
            I => \N__3664\
        );

    \I__770\ : LocalMux
    port map (
            O => \N__3708\,
            I => \N__3661\
        );

    \I__769\ : InMux
    port map (
            O => \N__3707\,
            I => \N__3656\
        );

    \I__768\ : InMux
    port map (
            O => \N__3706\,
            I => \N__3656\
        );

    \I__767\ : InMux
    port map (
            O => \N__3705\,
            I => \N__3649\
        );

    \I__766\ : InMux
    port map (
            O => \N__3704\,
            I => \N__3649\
        );

    \I__765\ : InMux
    port map (
            O => \N__3703\,
            I => \N__3649\
        );

    \I__764\ : InMux
    port map (
            O => \N__3700\,
            I => \N__3644\
        );

    \I__763\ : InMux
    port map (
            O => \N__3699\,
            I => \N__3644\
        );

    \I__762\ : InMux
    port map (
            O => \N__3698\,
            I => \N__3639\
        );

    \I__761\ : InMux
    port map (
            O => \N__3697\,
            I => \N__3639\
        );

    \I__760\ : Odrv4
    port map (
            O => \N__3694\,
            I => ctrl_tap_fsm_state_0
        );

    \I__759\ : LocalMux
    port map (
            O => \N__3689\,
            I => ctrl_tap_fsm_state_0
        );

    \I__758\ : LocalMux
    port map (
            O => \N__3680\,
            I => ctrl_tap_fsm_state_0
        );

    \I__757\ : LocalMux
    port map (
            O => \N__3677\,
            I => ctrl_tap_fsm_state_0
        );

    \I__756\ : LocalMux
    port map (
            O => \N__3672\,
            I => ctrl_tap_fsm_state_0
        );

    \I__755\ : LocalMux
    port map (
            O => \N__3669\,
            I => ctrl_tap_fsm_state_0
        );

    \I__754\ : LocalMux
    port map (
            O => \N__3664\,
            I => ctrl_tap_fsm_state_0
        );

    \I__753\ : Odrv4
    port map (
            O => \N__3661\,
            I => ctrl_tap_fsm_state_0
        );

    \I__752\ : LocalMux
    port map (
            O => \N__3656\,
            I => ctrl_tap_fsm_state_0
        );

    \I__751\ : LocalMux
    port map (
            O => \N__3649\,
            I => ctrl_tap_fsm_state_0
        );

    \I__750\ : LocalMux
    port map (
            O => \N__3644\,
            I => ctrl_tap_fsm_state_0
        );

    \I__749\ : LocalMux
    port map (
            O => \N__3639\,
            I => ctrl_tap_fsm_state_0
        );

    \I__748\ : CascadeMux
    port map (
            O => \N__3614\,
            I => \n17_cascade_\
        );

    \I__747\ : CascadeMux
    port map (
            O => \N__3611\,
            I => \n1687_cascade_\
        );

    \I__746\ : InMux
    port map (
            O => \N__3608\,
            I => \N__3605\
        );

    \I__745\ : LocalMux
    port map (
            O => \N__3605\,
            I => n2234
        );

    \I__744\ : InMux
    port map (
            O => \N__3602\,
            I => \N__3599\
        );

    \I__743\ : LocalMux
    port map (
            O => \N__3599\,
            I => n8
        );

    \I__742\ : InMux
    port map (
            O => \N__3596\,
            I => \N__3593\
        );

    \I__741\ : LocalMux
    port map (
            O => \N__3593\,
            I => n2198
        );

    \I__740\ : InMux
    port map (
            O => \N__3590\,
            I => \N__3586\
        );

    \I__739\ : InMux
    port map (
            O => \N__3589\,
            I => \N__3583\
        );

    \I__738\ : LocalMux
    port map (
            O => \N__3586\,
            I => \N__3580\
        );

    \I__737\ : LocalMux
    port map (
            O => \N__3583\,
            I => \ctrl_tap_instructionShift_0\
        );

    \I__736\ : Odrv12
    port map (
            O => \N__3580\,
            I => \ctrl_tap_instructionShift_0\
        );

    \I__735\ : InMux
    port map (
            O => \N__3575\,
            I => \N__3572\
        );

    \I__734\ : LocalMux
    port map (
            O => \N__3572\,
            I => ctrl_tap_bypass
        );

    \I__733\ : CascadeMux
    port map (
            O => \N__3569\,
            I => \n2198_cascade_\
        );

    \I__732\ : InMux
    port map (
            O => \N__3566\,
            I => \N__3563\
        );

    \I__731\ : LocalMux
    port map (
            O => \N__3563\,
            I => n4
        );

    \I__730\ : InMux
    port map (
            O => \N__3560\,
            I => \N__3557\
        );

    \I__729\ : LocalMux
    port map (
            O => \N__3557\,
            I => \ctrl_tap_tdoUnbufferd_N_213\
        );

    \I__728\ : CascadeMux
    port map (
            O => \N__3554\,
            I => \N__3551\
        );

    \I__727\ : InMux
    port map (
            O => \N__3551\,
            I => \N__3547\
        );

    \I__726\ : InMux
    port map (
            O => \N__3550\,
            I => \N__3544\
        );

    \I__725\ : LocalMux
    port map (
            O => \N__3547\,
            I => \ctrl_idcodeArea_shifter_27\
        );

    \I__724\ : LocalMux
    port map (
            O => \N__3544\,
            I => \ctrl_idcodeArea_shifter_27\
        );

    \I__723\ : CascadeMux
    port map (
            O => \N__3539\,
            I => \N__3535\
        );

    \I__722\ : CascadeMux
    port map (
            O => \N__3538\,
            I => \N__3532\
        );

    \I__721\ : InMux
    port map (
            O => \N__3535\,
            I => \N__3527\
        );

    \I__720\ : InMux
    port map (
            O => \N__3532\,
            I => \N__3527\
        );

    \I__719\ : LocalMux
    port map (
            O => \N__3527\,
            I => \ctrl_idcodeArea_shifter_26\
        );

    \I__718\ : InMux
    port map (
            O => \N__3524\,
            I => \N__3519\
        );

    \I__717\ : InMux
    port map (
            O => \N__3523\,
            I => \N__3516\
        );

    \I__716\ : InMux
    port map (
            O => \N__3522\,
            I => \N__3513\
        );

    \I__715\ : LocalMux
    port map (
            O => \N__3519\,
            I => \N__3509\
        );

    \I__714\ : LocalMux
    port map (
            O => \N__3516\,
            I => \N__3506\
        );

    \I__713\ : LocalMux
    port map (
            O => \N__3513\,
            I => \N__3503\
        );

    \I__712\ : InMux
    port map (
            O => \N__3512\,
            I => \N__3500\
        );

    \I__711\ : Span4Mux_v
    port map (
            O => \N__3509\,
            I => \N__3495\
        );

    \I__710\ : Span4Mux_h
    port map (
            O => \N__3506\,
            I => \N__3495\
        );

    \I__709\ : Span4Mux_v
    port map (
            O => \N__3503\,
            I => \N__3490\
        );

    \I__708\ : LocalMux
    port map (
            O => \N__3500\,
            I => \N__3490\
        );

    \I__707\ : Odrv4
    port map (
            O => \N__3495\,
            I => io_jtag_tdi_c
        );

    \I__706\ : Odrv4
    port map (
            O => \N__3490\,
            I => io_jtag_tdi_c
        );

    \I__705\ : CascadeMux
    port map (
            O => \N__3485\,
            I => \N__3481\
        );

    \I__704\ : InMux
    port map (
            O => \N__3484\,
            I => \N__3478\
        );

    \I__703\ : InMux
    port map (
            O => \N__3481\,
            I => \N__3475\
        );

    \I__702\ : LocalMux
    port map (
            O => \N__3478\,
            I => \ctrl_idcodeArea_shifter_23\
        );

    \I__701\ : LocalMux
    port map (
            O => \N__3475\,
            I => \ctrl_idcodeArea_shifter_23\
        );

    \I__700\ : CascadeMux
    port map (
            O => \N__3470\,
            I => \N__3466\
        );

    \I__699\ : InMux
    port map (
            O => \N__3469\,
            I => \N__3463\
        );

    \I__698\ : InMux
    port map (
            O => \N__3466\,
            I => \N__3460\
        );

    \I__697\ : LocalMux
    port map (
            O => \N__3463\,
            I => \ctrl_idcodeArea_shifter_22\
        );

    \I__696\ : LocalMux
    port map (
            O => \N__3460\,
            I => \ctrl_idcodeArea_shifter_22\
        );

    \I__695\ : InMux
    port map (
            O => \N__3455\,
            I => \N__3449\
        );

    \I__694\ : InMux
    port map (
            O => \N__3454\,
            I => \N__3449\
        );

    \I__693\ : LocalMux
    port map (
            O => \N__3449\,
            I => \ctrl_idcodeArea_shifter_21\
        );

    \I__692\ : CascadeMux
    port map (
            O => \N__3446\,
            I => \N__3442\
        );

    \I__691\ : InMux
    port map (
            O => \N__3445\,
            I => \N__3439\
        );

    \I__690\ : InMux
    port map (
            O => \N__3442\,
            I => \N__3436\
        );

    \I__689\ : LocalMux
    port map (
            O => \N__3439\,
            I => \ctrl_idcodeArea_shifter_18\
        );

    \I__688\ : LocalMux
    port map (
            O => \N__3436\,
            I => \ctrl_idcodeArea_shifter_18\
        );

    \I__687\ : CascadeMux
    port map (
            O => \N__3431\,
            I => \N__3397\
        );

    \I__686\ : InMux
    port map (
            O => \N__3430\,
            I => \N__3388\
        );

    \I__685\ : InMux
    port map (
            O => \N__3429\,
            I => \N__3388\
        );

    \I__684\ : InMux
    port map (
            O => \N__3428\,
            I => \N__3388\
        );

    \I__683\ : InMux
    port map (
            O => \N__3427\,
            I => \N__3388\
        );

    \I__682\ : InMux
    port map (
            O => \N__3426\,
            I => \N__3371\
        );

    \I__681\ : InMux
    port map (
            O => \N__3425\,
            I => \N__3371\
        );

    \I__680\ : InMux
    port map (
            O => \N__3424\,
            I => \N__3371\
        );

    \I__679\ : InMux
    port map (
            O => \N__3423\,
            I => \N__3371\
        );

    \I__678\ : InMux
    port map (
            O => \N__3422\,
            I => \N__3371\
        );

    \I__677\ : InMux
    port map (
            O => \N__3421\,
            I => \N__3371\
        );

    \I__676\ : InMux
    port map (
            O => \N__3420\,
            I => \N__3371\
        );

    \I__675\ : InMux
    port map (
            O => \N__3419\,
            I => \N__3371\
        );

    \I__674\ : InMux
    port map (
            O => \N__3418\,
            I => \N__3360\
        );

    \I__673\ : InMux
    port map (
            O => \N__3417\,
            I => \N__3360\
        );

    \I__672\ : InMux
    port map (
            O => \N__3416\,
            I => \N__3360\
        );

    \I__671\ : InMux
    port map (
            O => \N__3415\,
            I => \N__3360\
        );

    \I__670\ : InMux
    port map (
            O => \N__3414\,
            I => \N__3360\
        );

    \I__669\ : InMux
    port map (
            O => \N__3413\,
            I => \N__3349\
        );

    \I__668\ : InMux
    port map (
            O => \N__3412\,
            I => \N__3349\
        );

    \I__667\ : InMux
    port map (
            O => \N__3411\,
            I => \N__3349\
        );

    \I__666\ : InMux
    port map (
            O => \N__3410\,
            I => \N__3349\
        );

    \I__665\ : InMux
    port map (
            O => \N__3409\,
            I => \N__3349\
        );

    \I__664\ : InMux
    port map (
            O => \N__3408\,
            I => \N__3332\
        );

    \I__663\ : InMux
    port map (
            O => \N__3407\,
            I => \N__3332\
        );

    \I__662\ : InMux
    port map (
            O => \N__3406\,
            I => \N__3332\
        );

    \I__661\ : InMux
    port map (
            O => \N__3405\,
            I => \N__3332\
        );

    \I__660\ : InMux
    port map (
            O => \N__3404\,
            I => \N__3332\
        );

    \I__659\ : InMux
    port map (
            O => \N__3403\,
            I => \N__3332\
        );

    \I__658\ : InMux
    port map (
            O => \N__3402\,
            I => \N__3332\
        );

    \I__657\ : InMux
    port map (
            O => \N__3401\,
            I => \N__3332\
        );

    \I__656\ : InMux
    port map (
            O => \N__3400\,
            I => \N__3327\
        );

    \I__655\ : InMux
    port map (
            O => \N__3397\,
            I => \N__3327\
        );

    \I__654\ : LocalMux
    port map (
            O => \N__3388\,
            I => n15
        );

    \I__653\ : LocalMux
    port map (
            O => \N__3371\,
            I => n15
        );

    \I__652\ : LocalMux
    port map (
            O => \N__3360\,
            I => n15
        );

    \I__651\ : LocalMux
    port map (
            O => \N__3349\,
            I => n15
        );

    \I__650\ : LocalMux
    port map (
            O => \N__3332\,
            I => n15
        );

    \I__649\ : LocalMux
    port map (
            O => \N__3327\,
            I => n15
        );

    \I__648\ : CascadeMux
    port map (
            O => \N__3314\,
            I => \N__3310\
        );

    \I__647\ : CascadeMux
    port map (
            O => \N__3313\,
            I => \N__3307\
        );

    \I__646\ : InMux
    port map (
            O => \N__3310\,
            I => \N__3302\
        );

    \I__645\ : InMux
    port map (
            O => \N__3307\,
            I => \N__3302\
        );

    \I__644\ : LocalMux
    port map (
            O => \N__3302\,
            I => \ctrl_idcodeArea_shifter_20\
        );

    \I__643\ : CascadeMux
    port map (
            O => \N__3299\,
            I => \N__3287\
        );

    \I__642\ : CascadeMux
    port map (
            O => \N__3298\,
            I => \N__3282\
        );

    \I__641\ : CascadeMux
    port map (
            O => \N__3297\,
            I => \N__3279\
        );

    \I__640\ : CascadeMux
    port map (
            O => \N__3296\,
            I => \N__3275\
        );

    \I__639\ : CascadeMux
    port map (
            O => \N__3295\,
            I => \N__3272\
        );

    \I__638\ : CascadeMux
    port map (
            O => \N__3294\,
            I => \N__3267\
        );

    \I__637\ : CascadeMux
    port map (
            O => \N__3293\,
            I => \N__3263\
        );

    \I__636\ : CascadeMux
    port map (
            O => \N__3292\,
            I => \N__3260\
        );

    \I__635\ : InMux
    port map (
            O => \N__3291\,
            I => \N__3250\
        );

    \I__634\ : InMux
    port map (
            O => \N__3290\,
            I => \N__3250\
        );

    \I__633\ : InMux
    port map (
            O => \N__3287\,
            I => \N__3250\
        );

    \I__632\ : InMux
    port map (
            O => \N__3286\,
            I => \N__3250\
        );

    \I__631\ : InMux
    port map (
            O => \N__3285\,
            I => \N__3220\
        );

    \I__630\ : InMux
    port map (
            O => \N__3282\,
            I => \N__3220\
        );

    \I__629\ : InMux
    port map (
            O => \N__3279\,
            I => \N__3220\
        );

    \I__628\ : InMux
    port map (
            O => \N__3278\,
            I => \N__3220\
        );

    \I__627\ : InMux
    port map (
            O => \N__3275\,
            I => \N__3220\
        );

    \I__626\ : InMux
    port map (
            O => \N__3272\,
            I => \N__3220\
        );

    \I__625\ : InMux
    port map (
            O => \N__3271\,
            I => \N__3220\
        );

    \I__624\ : InMux
    port map (
            O => \N__3270\,
            I => \N__3220\
        );

    \I__623\ : InMux
    port map (
            O => \N__3267\,
            I => \N__3209\
        );

    \I__622\ : InMux
    port map (
            O => \N__3266\,
            I => \N__3209\
        );

    \I__621\ : InMux
    port map (
            O => \N__3263\,
            I => \N__3209\
        );

    \I__620\ : InMux
    port map (
            O => \N__3260\,
            I => \N__3209\
        );

    \I__619\ : InMux
    port map (
            O => \N__3259\,
            I => \N__3209\
        );

    \I__618\ : LocalMux
    port map (
            O => \N__3250\,
            I => \N__3200\
        );

    \I__617\ : InMux
    port map (
            O => \N__3249\,
            I => \N__3193\
        );

    \I__616\ : InMux
    port map (
            O => \N__3248\,
            I => \N__3193\
        );

    \I__615\ : InMux
    port map (
            O => \N__3247\,
            I => \N__3193\
        );

    \I__614\ : InMux
    port map (
            O => \N__3246\,
            I => \N__3188\
        );

    \I__613\ : InMux
    port map (
            O => \N__3245\,
            I => \N__3188\
        );

    \I__612\ : InMux
    port map (
            O => \N__3244\,
            I => \N__3179\
        );

    \I__611\ : InMux
    port map (
            O => \N__3243\,
            I => \N__3179\
        );

    \I__610\ : InMux
    port map (
            O => \N__3242\,
            I => \N__3179\
        );

    \I__609\ : InMux
    port map (
            O => \N__3241\,
            I => \N__3179\
        );

    \I__608\ : InMux
    port map (
            O => \N__3240\,
            I => \N__3170\
        );

    \I__607\ : InMux
    port map (
            O => \N__3239\,
            I => \N__3170\
        );

    \I__606\ : InMux
    port map (
            O => \N__3238\,
            I => \N__3170\
        );

    \I__605\ : InMux
    port map (
            O => \N__3237\,
            I => \N__3170\
        );

    \I__604\ : LocalMux
    port map (
            O => \N__3220\,
            I => \N__3165\
        );

    \I__603\ : LocalMux
    port map (
            O => \N__3209\,
            I => \N__3165\
        );

    \I__602\ : InMux
    port map (
            O => \N__3208\,
            I => \N__3160\
        );

    \I__601\ : InMux
    port map (
            O => \N__3207\,
            I => \N__3160\
        );

    \I__600\ : InMux
    port map (
            O => \N__3206\,
            I => \N__3151\
        );

    \I__599\ : InMux
    port map (
            O => \N__3205\,
            I => \N__3151\
        );

    \I__598\ : InMux
    port map (
            O => \N__3204\,
            I => \N__3151\
        );

    \I__597\ : InMux
    port map (
            O => \N__3203\,
            I => \N__3151\
        );

    \I__596\ : Odrv4
    port map (
            O => \N__3200\,
            I => n1489
        );

    \I__595\ : LocalMux
    port map (
            O => \N__3193\,
            I => n1489
        );

    \I__594\ : LocalMux
    port map (
            O => \N__3188\,
            I => n1489
        );

    \I__593\ : LocalMux
    port map (
            O => \N__3179\,
            I => n1489
        );

    \I__592\ : LocalMux
    port map (
            O => \N__3170\,
            I => n1489
        );

    \I__591\ : Odrv4
    port map (
            O => \N__3165\,
            I => n1489
        );

    \I__590\ : LocalMux
    port map (
            O => \N__3160\,
            I => n1489
        );

    \I__589\ : LocalMux
    port map (
            O => \N__3151\,
            I => n1489
        );

    \I__588\ : CascadeMux
    port map (
            O => \N__3134\,
            I => \N__3130\
        );

    \I__587\ : InMux
    port map (
            O => \N__3133\,
            I => \N__3125\
        );

    \I__586\ : InMux
    port map (
            O => \N__3130\,
            I => \N__3125\
        );

    \I__585\ : LocalMux
    port map (
            O => \N__3125\,
            I => \ctrl_idcodeArea_shifter_19\
        );

    \I__584\ : CascadeMux
    port map (
            O => \N__3122\,
            I => \n2185_cascade_\
        );

    \I__583\ : InMux
    port map (
            O => \N__3119\,
            I => \N__3099\
        );

    \I__582\ : InMux
    port map (
            O => \N__3118\,
            I => \N__3099\
        );

    \I__581\ : InMux
    port map (
            O => \N__3117\,
            I => \N__3099\
        );

    \I__580\ : InMux
    port map (
            O => \N__3116\,
            I => \N__3099\
        );

    \I__579\ : InMux
    port map (
            O => \N__3115\,
            I => \N__3079\
        );

    \I__578\ : InMux
    port map (
            O => \N__3114\,
            I => \N__3079\
        );

    \I__577\ : InMux
    port map (
            O => \N__3113\,
            I => \N__3079\
        );

    \I__576\ : InMux
    port map (
            O => \N__3112\,
            I => \N__3079\
        );

    \I__575\ : InMux
    port map (
            O => \N__3111\,
            I => \N__3070\
        );

    \I__574\ : InMux
    port map (
            O => \N__3110\,
            I => \N__3070\
        );

    \I__573\ : InMux
    port map (
            O => \N__3109\,
            I => \N__3070\
        );

    \I__572\ : InMux
    port map (
            O => \N__3108\,
            I => \N__3070\
        );

    \I__571\ : LocalMux
    port map (
            O => \N__3099\,
            I => \N__3067\
        );

    \I__570\ : InMux
    port map (
            O => \N__3098\,
            I => \N__3058\
        );

    \I__569\ : InMux
    port map (
            O => \N__3097\,
            I => \N__3058\
        );

    \I__568\ : InMux
    port map (
            O => \N__3096\,
            I => \N__3058\
        );

    \I__567\ : InMux
    port map (
            O => \N__3095\,
            I => \N__3058\
        );

    \I__566\ : InMux
    port map (
            O => \N__3094\,
            I => \N__3051\
        );

    \I__565\ : InMux
    port map (
            O => \N__3093\,
            I => \N__3051\
        );

    \I__564\ : InMux
    port map (
            O => \N__3092\,
            I => \N__3051\
        );

    \I__563\ : InMux
    port map (
            O => \N__3091\,
            I => \N__3042\
        );

    \I__562\ : InMux
    port map (
            O => \N__3090\,
            I => \N__3042\
        );

    \I__561\ : InMux
    port map (
            O => \N__3089\,
            I => \N__3042\
        );

    \I__560\ : InMux
    port map (
            O => \N__3088\,
            I => \N__3042\
        );

    \I__559\ : LocalMux
    port map (
            O => \N__3079\,
            I => n1848
        );

    \I__558\ : LocalMux
    port map (
            O => \N__3070\,
            I => n1848
        );

    \I__557\ : Odrv4
    port map (
            O => \N__3067\,
            I => n1848
        );

    \I__556\ : LocalMux
    port map (
            O => \N__3058\,
            I => n1848
        );

    \I__555\ : LocalMux
    port map (
            O => \N__3051\,
            I => n1848
        );

    \I__554\ : LocalMux
    port map (
            O => \N__3042\,
            I => n1848
        );

    \I__553\ : InMux
    port map (
            O => \N__3029\,
            I => \N__3025\
        );

    \I__552\ : InMux
    port map (
            O => \N__3028\,
            I => \N__3022\
        );

    \I__551\ : LocalMux
    port map (
            O => \N__3025\,
            I => \myClockArea_timeout_counter_value_7\
        );

    \I__550\ : LocalMux
    port map (
            O => \N__3022\,
            I => \myClockArea_timeout_counter_value_7\
        );

    \I__549\ : InMux
    port map (
            O => \N__3017\,
            I => \N__3013\
        );

    \I__548\ : InMux
    port map (
            O => \N__3016\,
            I => \N__3010\
        );

    \I__547\ : LocalMux
    port map (
            O => \N__3013\,
            I => \myClockArea_timeout_counter_value_21\
        );

    \I__546\ : LocalMux
    port map (
            O => \N__3010\,
            I => \myClockArea_timeout_counter_value_21\
        );

    \I__545\ : InMux
    port map (
            O => \N__3005\,
            I => \N__3002\
        );

    \I__544\ : LocalMux
    port map (
            O => \N__3002\,
            I => n11
        );

    \I__543\ : InMux
    port map (
            O => \N__2999\,
            I => \N__2995\
        );

    \I__542\ : InMux
    port map (
            O => \N__2998\,
            I => \N__2992\
        );

    \I__541\ : LocalMux
    port map (
            O => \N__2995\,
            I => \myClockArea_timeout_counter_value_19\
        );

    \I__540\ : LocalMux
    port map (
            O => \N__2992\,
            I => \myClockArea_timeout_counter_value_19\
        );

    \I__539\ : InMux
    port map (
            O => \N__2987\,
            I => \N__2983\
        );

    \I__538\ : InMux
    port map (
            O => \N__2986\,
            I => \N__2980\
        );

    \I__537\ : LocalMux
    port map (
            O => \N__2983\,
            I => \myClockArea_timeout_counter_value_15\
        );

    \I__536\ : LocalMux
    port map (
            O => \N__2980\,
            I => \myClockArea_timeout_counter_value_15\
        );

    \I__535\ : CascadeMux
    port map (
            O => \N__2975\,
            I => \N__2971\
        );

    \I__534\ : InMux
    port map (
            O => \N__2974\,
            I => \N__2968\
        );

    \I__533\ : InMux
    port map (
            O => \N__2971\,
            I => \N__2965\
        );

    \I__532\ : LocalMux
    port map (
            O => \N__2968\,
            I => \myClockArea_timeout_counter_value_20\
        );

    \I__531\ : LocalMux
    port map (
            O => \N__2965\,
            I => \myClockArea_timeout_counter_value_20\
        );

    \I__530\ : InMux
    port map (
            O => \N__2960\,
            I => \N__2956\
        );

    \I__529\ : InMux
    port map (
            O => \N__2959\,
            I => \N__2953\
        );

    \I__528\ : LocalMux
    port map (
            O => \N__2956\,
            I => \myClockArea_timeout_counter_value_11\
        );

    \I__527\ : LocalMux
    port map (
            O => \N__2953\,
            I => \myClockArea_timeout_counter_value_11\
        );

    \I__526\ : InMux
    port map (
            O => \N__2948\,
            I => \N__2945\
        );

    \I__525\ : LocalMux
    port map (
            O => \N__2945\,
            I => n2220
        );

    \I__524\ : InMux
    port map (
            O => \N__2942\,
            I => \N__2938\
        );

    \I__523\ : InMux
    port map (
            O => \N__2941\,
            I => \N__2935\
        );

    \I__522\ : LocalMux
    port map (
            O => \N__2938\,
            I => \myClockArea_timeout_counter_value_9\
        );

    \I__521\ : LocalMux
    port map (
            O => \N__2935\,
            I => \myClockArea_timeout_counter_value_9\
        );

    \I__520\ : InMux
    port map (
            O => \N__2930\,
            I => \N__2926\
        );

    \I__519\ : InMux
    port map (
            O => \N__2929\,
            I => \N__2923\
        );

    \I__518\ : LocalMux
    port map (
            O => \N__2926\,
            I => \myClockArea_timeout_counter_value_18\
        );

    \I__517\ : LocalMux
    port map (
            O => \N__2923\,
            I => \myClockArea_timeout_counter_value_18\
        );

    \I__516\ : CascadeMux
    port map (
            O => \N__2918\,
            I => \N__2914\
        );

    \I__515\ : InMux
    port map (
            O => \N__2917\,
            I => \N__2911\
        );

    \I__514\ : InMux
    port map (
            O => \N__2914\,
            I => \N__2908\
        );

    \I__513\ : LocalMux
    port map (
            O => \N__2911\,
            I => \myClockArea_timeout_counter_value_12\
        );

    \I__512\ : LocalMux
    port map (
            O => \N__2908\,
            I => \myClockArea_timeout_counter_value_12\
        );

    \I__511\ : InMux
    port map (
            O => \N__2903\,
            I => \N__2899\
        );

    \I__510\ : InMux
    port map (
            O => \N__2902\,
            I => \N__2896\
        );

    \I__509\ : LocalMux
    port map (
            O => \N__2899\,
            I => \myClockArea_timeout_counter_value_14\
        );

    \I__508\ : LocalMux
    port map (
            O => \N__2896\,
            I => \myClockArea_timeout_counter_value_14\
        );

    \I__507\ : InMux
    port map (
            O => \N__2891\,
            I => \N__2888\
        );

    \I__506\ : LocalMux
    port map (
            O => \N__2888\,
            I => n13
        );

    \I__505\ : InMux
    port map (
            O => \N__2885\,
            I => \N__2880\
        );

    \I__504\ : InMux
    port map (
            O => \N__2884\,
            I => \N__2877\
        );

    \I__503\ : InMux
    port map (
            O => \N__2883\,
            I => \N__2874\
        );

    \I__502\ : LocalMux
    port map (
            O => \N__2880\,
            I => \N__2871\
        );

    \I__501\ : LocalMux
    port map (
            O => \N__2877\,
            I => \myClockArea_timeout_state\
        );

    \I__500\ : LocalMux
    port map (
            O => \N__2874\,
            I => \myClockArea_timeout_state\
        );

    \I__499\ : Odrv4
    port map (
            O => \N__2871\,
            I => \myClockArea_timeout_state\
        );

    \I__498\ : IoInMux
    port map (
            O => \N__2864\,
            I => \N__2861\
        );

    \I__497\ : LocalMux
    port map (
            O => \N__2861\,
            I => \N__2857\
        );

    \I__496\ : InMux
    port map (
            O => \N__2860\,
            I => \N__2854\
        );

    \I__495\ : Odrv12
    port map (
            O => \N__2857\,
            I => io_leds_c_3
        );

    \I__494\ : LocalMux
    port map (
            O => \N__2854\,
            I => io_leds_c_3
        );

    \I__493\ : ClkMux
    port map (
            O => \N__2849\,
            I => \N__2834\
        );

    \I__492\ : ClkMux
    port map (
            O => \N__2848\,
            I => \N__2834\
        );

    \I__491\ : ClkMux
    port map (
            O => \N__2847\,
            I => \N__2834\
        );

    \I__490\ : ClkMux
    port map (
            O => \N__2846\,
            I => \N__2834\
        );

    \I__489\ : ClkMux
    port map (
            O => \N__2845\,
            I => \N__2834\
        );

    \I__488\ : GlobalMux
    port map (
            O => \N__2834\,
            I => \N__2831\
        );

    \I__487\ : gio2CtrlBuf
    port map (
            O => \N__2831\,
            I => global_clk_c
        );

    \I__486\ : InMux
    port map (
            O => \N__2828\,
            I => \N__2822\
        );

    \I__485\ : InMux
    port map (
            O => \N__2827\,
            I => \N__2822\
        );

    \I__484\ : LocalMux
    port map (
            O => \N__2822\,
            I => \ctrl_idcodeArea_shifter_25\
        );

    \I__483\ : CascadeMux
    port map (
            O => \N__2819\,
            I => \N__2815\
        );

    \I__482\ : InMux
    port map (
            O => \N__2818\,
            I => \N__2810\
        );

    \I__481\ : InMux
    port map (
            O => \N__2815\,
            I => \N__2810\
        );

    \I__480\ : LocalMux
    port map (
            O => \N__2810\,
            I => \ctrl_idcodeArea_shifter_24\
        );

    \I__479\ : IoInMux
    port map (
            O => \N__2807\,
            I => \N__2804\
        );

    \I__478\ : LocalMux
    port map (
            O => \N__2804\,
            I => \N__2801\
        );

    \I__477\ : IoSpan4Mux
    port map (
            O => \N__2801\,
            I => \N__2797\
        );

    \I__476\ : CascadeMux
    port map (
            O => \N__2800\,
            I => \N__2793\
        );

    \I__475\ : Span4Mux_s3_h
    port map (
            O => \N__2797\,
            I => \N__2790\
        );

    \I__474\ : InMux
    port map (
            O => \N__2796\,
            I => \N__2787\
        );

    \I__473\ : InMux
    port map (
            O => \N__2793\,
            I => \N__2784\
        );

    \I__472\ : Odrv4
    port map (
            O => \N__2790\,
            I => io_leds_c_7
        );

    \I__471\ : LocalMux
    port map (
            O => \N__2787\,
            I => io_leds_c_7
        );

    \I__470\ : LocalMux
    port map (
            O => \N__2784\,
            I => io_leds_c_7
        );

    \I__469\ : InMux
    port map (
            O => \N__2777\,
            I => \N__2773\
        );

    \I__468\ : InMux
    port map (
            O => \N__2776\,
            I => \N__2770\
        );

    \I__467\ : LocalMux
    port map (
            O => \N__2773\,
            I => \myClockArea_timeout_counter_value_3\
        );

    \I__466\ : LocalMux
    port map (
            O => \N__2770\,
            I => \myClockArea_timeout_counter_value_3\
        );

    \I__465\ : InMux
    port map (
            O => \N__2765\,
            I => \N__2761\
        );

    \I__464\ : InMux
    port map (
            O => \N__2764\,
            I => \N__2758\
        );

    \I__463\ : LocalMux
    port map (
            O => \N__2761\,
            I => \myClockArea_timeout_counter_value_1\
        );

    \I__462\ : LocalMux
    port map (
            O => \N__2758\,
            I => \myClockArea_timeout_counter_value_1\
        );

    \I__461\ : CascadeMux
    port map (
            O => \N__2753\,
            I => \N__2749\
        );

    \I__460\ : InMux
    port map (
            O => \N__2752\,
            I => \N__2746\
        );

    \I__459\ : InMux
    port map (
            O => \N__2749\,
            I => \N__2743\
        );

    \I__458\ : LocalMux
    port map (
            O => \N__2746\,
            I => \myClockArea_timeout_counter_value_5\
        );

    \I__457\ : LocalMux
    port map (
            O => \N__2743\,
            I => \myClockArea_timeout_counter_value_5\
        );

    \I__456\ : InMux
    port map (
            O => \N__2738\,
            I => \N__2734\
        );

    \I__455\ : InMux
    port map (
            O => \N__2737\,
            I => \N__2731\
        );

    \I__454\ : LocalMux
    port map (
            O => \N__2734\,
            I => \myClockArea_timeout_counter_value_0\
        );

    \I__453\ : LocalMux
    port map (
            O => \N__2731\,
            I => \myClockArea_timeout_counter_value_0\
        );

    \I__452\ : InMux
    port map (
            O => \N__2726\,
            I => \N__2723\
        );

    \I__451\ : LocalMux
    port map (
            O => \N__2723\,
            I => n2309
        );

    \I__450\ : InMux
    port map (
            O => \N__2720\,
            I => \N__2716\
        );

    \I__449\ : InMux
    port map (
            O => \N__2719\,
            I => \N__2713\
        );

    \I__448\ : LocalMux
    port map (
            O => \N__2716\,
            I => \myClockArea_timeout_counter_value_4\
        );

    \I__447\ : LocalMux
    port map (
            O => \N__2713\,
            I => \myClockArea_timeout_counter_value_4\
        );

    \I__446\ : InMux
    port map (
            O => \N__2708\,
            I => \N__2704\
        );

    \I__445\ : InMux
    port map (
            O => \N__2707\,
            I => \N__2701\
        );

    \I__444\ : LocalMux
    port map (
            O => \N__2704\,
            I => \myClockArea_timeout_counter_value_6\
        );

    \I__443\ : LocalMux
    port map (
            O => \N__2701\,
            I => \myClockArea_timeout_counter_value_6\
        );

    \I__442\ : CascadeMux
    port map (
            O => \N__2696\,
            I => \N__2692\
        );

    \I__441\ : InMux
    port map (
            O => \N__2695\,
            I => \N__2689\
        );

    \I__440\ : InMux
    port map (
            O => \N__2692\,
            I => \N__2686\
        );

    \I__439\ : LocalMux
    port map (
            O => \N__2689\,
            I => \myClockArea_timeout_counter_value_22\
        );

    \I__438\ : LocalMux
    port map (
            O => \N__2686\,
            I => \myClockArea_timeout_counter_value_22\
        );

    \I__437\ : InMux
    port map (
            O => \N__2681\,
            I => \N__2677\
        );

    \I__436\ : InMux
    port map (
            O => \N__2680\,
            I => \N__2674\
        );

    \I__435\ : LocalMux
    port map (
            O => \N__2677\,
            I => \myClockArea_timeout_counter_value_16\
        );

    \I__434\ : LocalMux
    port map (
            O => \N__2674\,
            I => \myClockArea_timeout_counter_value_16\
        );

    \I__433\ : InMux
    port map (
            O => \N__2669\,
            I => \N__2665\
        );

    \I__432\ : InMux
    port map (
            O => \N__2668\,
            I => \N__2662\
        );

    \I__431\ : LocalMux
    port map (
            O => \N__2665\,
            I => \myClockArea_timeout_counter_value_17\
        );

    \I__430\ : LocalMux
    port map (
            O => \N__2662\,
            I => \myClockArea_timeout_counter_value_17\
        );

    \I__429\ : InMux
    port map (
            O => \N__2657\,
            I => \N__2653\
        );

    \I__428\ : InMux
    port map (
            O => \N__2656\,
            I => \N__2650\
        );

    \I__427\ : LocalMux
    port map (
            O => \N__2653\,
            I => \myClockArea_timeout_counter_value_8\
        );

    \I__426\ : LocalMux
    port map (
            O => \N__2650\,
            I => \myClockArea_timeout_counter_value_8\
        );

    \I__425\ : CascadeMux
    port map (
            O => \N__2645\,
            I => \N__2641\
        );

    \I__424\ : InMux
    port map (
            O => \N__2644\,
            I => \N__2638\
        );

    \I__423\ : InMux
    port map (
            O => \N__2641\,
            I => \N__2635\
        );

    \I__422\ : LocalMux
    port map (
            O => \N__2638\,
            I => \myClockArea_timeout_counter_value_10\
        );

    \I__421\ : LocalMux
    port map (
            O => \N__2635\,
            I => \myClockArea_timeout_counter_value_10\
        );

    \I__420\ : InMux
    port map (
            O => \N__2630\,
            I => \N__2626\
        );

    \I__419\ : InMux
    port map (
            O => \N__2629\,
            I => \N__2623\
        );

    \I__418\ : LocalMux
    port map (
            O => \N__2626\,
            I => \myClockArea_timeout_counter_value_2\
        );

    \I__417\ : LocalMux
    port map (
            O => \N__2623\,
            I => \myClockArea_timeout_counter_value_2\
        );

    \I__416\ : InMux
    port map (
            O => \N__2618\,
            I => \N__2615\
        );

    \I__415\ : LocalMux
    port map (
            O => \N__2615\,
            I => n2216
        );

    \I__414\ : CascadeMux
    port map (
            O => \N__2612\,
            I => \n2218_cascade_\
        );

    \I__413\ : InMux
    port map (
            O => \N__2609\,
            I => \N__2606\
        );

    \I__412\ : LocalMux
    port map (
            O => \N__2606\,
            I => n2222
        );

    \I__411\ : InMux
    port map (
            O => \N__2603\,
            I => \N__2599\
        );

    \I__410\ : InMux
    port map (
            O => \N__2602\,
            I => \N__2596\
        );

    \I__409\ : LocalMux
    port map (
            O => \N__2599\,
            I => \myClockArea_timeout_counter_value_13\
        );

    \I__408\ : LocalMux
    port map (
            O => \N__2596\,
            I => \myClockArea_timeout_counter_value_13\
        );

    \I__407\ : CascadeMux
    port map (
            O => \N__2591\,
            I => \n2228_cascade_\
        );

    \I__406\ : InMux
    port map (
            O => \N__2588\,
            I => \N__2585\
        );

    \I__405\ : LocalMux
    port map (
            O => \N__2585\,
            I => \N__2582\
        );

    \I__404\ : Odrv4
    port map (
            O => \N__2582\,
            I => n2185
        );

    \I__403\ : CascadeMux
    port map (
            O => \N__2579\,
            I => \n2282_cascade_\
        );

    \I__402\ : CascadeMux
    port map (
            O => \N__2576\,
            I => \n2326_cascade_\
        );

    \I__401\ : InMux
    port map (
            O => \N__2573\,
            I => \N__2570\
        );

    \I__400\ : LocalMux
    port map (
            O => \N__2570\,
            I => n2306
        );

    \I__399\ : CascadeMux
    port map (
            O => \N__2567\,
            I => \N__2563\
        );

    \I__398\ : CEMux
    port map (
            O => \N__2566\,
            I => \N__2560\
        );

    \I__397\ : InMux
    port map (
            O => \N__2563\,
            I => \N__2557\
        );

    \I__396\ : LocalMux
    port map (
            O => \N__2560\,
            I => n1022
        );

    \I__395\ : LocalMux
    port map (
            O => \N__2557\,
            I => n1022
        );

    \I__394\ : CascadeMux
    port map (
            O => \N__2552\,
            I => \n2231_cascade_\
        );

    \I__393\ : InMux
    port map (
            O => \N__2549\,
            I => \N__2546\
        );

    \I__392\ : LocalMux
    port map (
            O => \N__2546\,
            I => n2273
        );

    \I__391\ : CascadeMux
    port map (
            O => \N__2543\,
            I => \n2263_cascade_\
        );

    \I__390\ : InMux
    port map (
            O => \N__2540\,
            I => \N__2537\
        );

    \I__389\ : LocalMux
    port map (
            O => \N__2537\,
            I => n2323
        );

    \I__388\ : InMux
    port map (
            O => \N__2534\,
            I => \N__2531\
        );

    \I__387\ : LocalMux
    port map (
            O => \N__2531\,
            I => n2272
        );

    \I__386\ : CascadeMux
    port map (
            O => \N__2528\,
            I => \n1489_cascade_\
        );

    \I__385\ : CascadeMux
    port map (
            O => \N__2525\,
            I => \n1269_cascade_\
        );

    \I__384\ : InMux
    port map (
            O => \N__2522\,
            I => \N__2515\
        );

    \I__383\ : InMux
    port map (
            O => \N__2521\,
            I => \N__2512\
        );

    \I__382\ : InMux
    port map (
            O => \N__2520\,
            I => \N__2509\
        );

    \I__381\ : InMux
    port map (
            O => \N__2519\,
            I => \N__2504\
        );

    \I__380\ : InMux
    port map (
            O => \N__2518\,
            I => \N__2504\
        );

    \I__379\ : LocalMux
    port map (
            O => \N__2515\,
            I => ctrl_tap_instruction_0
        );

    \I__378\ : LocalMux
    port map (
            O => \N__2512\,
            I => ctrl_tap_instruction_0
        );

    \I__377\ : LocalMux
    port map (
            O => \N__2509\,
            I => ctrl_tap_instruction_0
        );

    \I__376\ : LocalMux
    port map (
            O => \N__2504\,
            I => ctrl_tap_instruction_0
        );

    \I__375\ : CascadeMux
    port map (
            O => \N__2495\,
            I => \N__2492\
        );

    \I__374\ : InMux
    port map (
            O => \N__2492\,
            I => \N__2488\
        );

    \I__373\ : InMux
    port map (
            O => \N__2491\,
            I => \N__2485\
        );

    \I__372\ : LocalMux
    port map (
            O => \N__2488\,
            I => \ctrl_tap_instructionShift_3\
        );

    \I__371\ : LocalMux
    port map (
            O => \N__2485\,
            I => \ctrl_tap_instructionShift_3\
        );

    \I__370\ : InMux
    port map (
            O => \N__2480\,
            I => \N__2476\
        );

    \I__369\ : CascadeMux
    port map (
            O => \N__2479\,
            I => \N__2471\
        );

    \I__368\ : LocalMux
    port map (
            O => \N__2476\,
            I => \N__2467\
        );

    \I__367\ : InMux
    port map (
            O => \N__2475\,
            I => \N__2464\
        );

    \I__366\ : InMux
    port map (
            O => \N__2474\,
            I => \N__2461\
        );

    \I__365\ : InMux
    port map (
            O => \N__2471\,
            I => \N__2456\
        );

    \I__364\ : InMux
    port map (
            O => \N__2470\,
            I => \N__2456\
        );

    \I__363\ : Odrv4
    port map (
            O => \N__2467\,
            I => ctrl_tap_instruction_3
        );

    \I__362\ : LocalMux
    port map (
            O => \N__2464\,
            I => ctrl_tap_instruction_3
        );

    \I__361\ : LocalMux
    port map (
            O => \N__2461\,
            I => ctrl_tap_instruction_3
        );

    \I__360\ : LocalMux
    port map (
            O => \N__2456\,
            I => ctrl_tap_instruction_3
        );

    \I__359\ : CascadeMux
    port map (
            O => \N__2447\,
            I => \N__2444\
        );

    \I__358\ : InMux
    port map (
            O => \N__2444\,
            I => \N__2440\
        );

    \I__357\ : InMux
    port map (
            O => \N__2443\,
            I => \N__2437\
        );

    \I__356\ : LocalMux
    port map (
            O => \N__2440\,
            I => \ctrl_tap_instructionShift_2\
        );

    \I__355\ : LocalMux
    port map (
            O => \N__2437\,
            I => \ctrl_tap_instructionShift_2\
        );

    \I__354\ : InMux
    port map (
            O => \N__2432\,
            I => \N__2425\
        );

    \I__353\ : InMux
    port map (
            O => \N__2431\,
            I => \N__2422\
        );

    \I__352\ : InMux
    port map (
            O => \N__2430\,
            I => \N__2419\
        );

    \I__351\ : InMux
    port map (
            O => \N__2429\,
            I => \N__2414\
        );

    \I__350\ : InMux
    port map (
            O => \N__2428\,
            I => \N__2414\
        );

    \I__349\ : LocalMux
    port map (
            O => \N__2425\,
            I => ctrl_tap_instruction_2
        );

    \I__348\ : LocalMux
    port map (
            O => \N__2422\,
            I => ctrl_tap_instruction_2
        );

    \I__347\ : LocalMux
    port map (
            O => \N__2419\,
            I => ctrl_tap_instruction_2
        );

    \I__346\ : LocalMux
    port map (
            O => \N__2414\,
            I => ctrl_tap_instruction_2
        );

    \I__345\ : InMux
    port map (
            O => \N__2405\,
            I => \N__2396\
        );

    \I__344\ : InMux
    port map (
            O => \N__2404\,
            I => \N__2396\
        );

    \I__343\ : InMux
    port map (
            O => \N__2403\,
            I => \N__2396\
        );

    \I__342\ : LocalMux
    port map (
            O => \N__2396\,
            I => n1269
        );

    \I__341\ : CascadeMux
    port map (
            O => \N__2393\,
            I => \N__2390\
        );

    \I__340\ : InMux
    port map (
            O => \N__2390\,
            I => \N__2386\
        );

    \I__339\ : InMux
    port map (
            O => \N__2389\,
            I => \N__2383\
        );

    \I__338\ : LocalMux
    port map (
            O => \N__2386\,
            I => \ctrl_tap_instructionShift_1\
        );

    \I__337\ : LocalMux
    port map (
            O => \N__2383\,
            I => \ctrl_tap_instructionShift_1\
        );

    \I__336\ : CascadeMux
    port map (
            O => \N__2378\,
            I => \N__2373\
        );

    \I__335\ : InMux
    port map (
            O => \N__2377\,
            I => \N__2368\
        );

    \I__334\ : InMux
    port map (
            O => \N__2376\,
            I => \N__2365\
        );

    \I__333\ : InMux
    port map (
            O => \N__2373\,
            I => \N__2362\
        );

    \I__332\ : InMux
    port map (
            O => \N__2372\,
            I => \N__2359\
        );

    \I__331\ : InMux
    port map (
            O => \N__2371\,
            I => \N__2356\
        );

    \I__330\ : LocalMux
    port map (
            O => \N__2368\,
            I => ctrl_tap_instruction_1
        );

    \I__329\ : LocalMux
    port map (
            O => \N__2365\,
            I => ctrl_tap_instruction_1
        );

    \I__328\ : LocalMux
    port map (
            O => \N__2362\,
            I => ctrl_tap_instruction_1
        );

    \I__327\ : LocalMux
    port map (
            O => \N__2359\,
            I => ctrl_tap_instruction_1
        );

    \I__326\ : LocalMux
    port map (
            O => \N__2356\,
            I => ctrl_tap_instruction_1
        );

    \I__325\ : InMux
    port map (
            O => \N__2345\,
            I => \N__2342\
        );

    \I__324\ : LocalMux
    port map (
            O => \N__2342\,
            I => n2248
        );

    \I__323\ : CascadeMux
    port map (
            O => \N__2339\,
            I => \n118_cascade_\
        );

    \I__322\ : CascadeMux
    port map (
            O => \N__2336\,
            I => \N__2333\
        );

    \I__321\ : InMux
    port map (
            O => \N__2333\,
            I => \N__2329\
        );

    \I__320\ : InMux
    port map (
            O => \N__2332\,
            I => \N__2326\
        );

    \I__319\ : LocalMux
    port map (
            O => \N__2329\,
            I => \N__2323\
        );

    \I__318\ : LocalMux
    port map (
            O => \N__2326\,
            I => \ctrl_idcodeArea_shifter_17\
        );

    \I__317\ : Odrv12
    port map (
            O => \N__2323\,
            I => \ctrl_idcodeArea_shifter_17\
        );

    \I__316\ : InMux
    port map (
            O => \N__2318\,
            I => \N__2314\
        );

    \I__315\ : InMux
    port map (
            O => \N__2317\,
            I => \N__2311\
        );

    \I__314\ : LocalMux
    port map (
            O => \N__2314\,
            I => \ctrl_idcodeArea_shifter_1\
        );

    \I__313\ : LocalMux
    port map (
            O => \N__2311\,
            I => \ctrl_idcodeArea_shifter_1\
        );

    \I__312\ : CascadeMux
    port map (
            O => \N__2306\,
            I => \n6_cascade_\
        );

    \I__311\ : InMux
    port map (
            O => \N__2303\,
            I => \N__2297\
        );

    \I__310\ : InMux
    port map (
            O => \N__2302\,
            I => \N__2297\
        );

    \I__309\ : LocalMux
    port map (
            O => \N__2297\,
            I => \ctrl_idcodeArea_shifter_0\
        );

    \I__308\ : InMux
    port map (
            O => \N__2294\,
            I => \N__2291\
        );

    \I__307\ : LocalMux
    port map (
            O => \N__2291\,
            I => n2085
        );

    \I__306\ : CascadeMux
    port map (
            O => \N__2288\,
            I => \n15_cascade_\
        );

    \I__305\ : CascadeMux
    port map (
            O => \N__2285\,
            I => \N__2281\
        );

    \I__304\ : InMux
    port map (
            O => \N__2284\,
            I => \N__2278\
        );

    \I__303\ : InMux
    port map (
            O => \N__2281\,
            I => \N__2275\
        );

    \I__302\ : LocalMux
    port map (
            O => \N__2278\,
            I => \N__2272\
        );

    \I__301\ : LocalMux
    port map (
            O => \N__2275\,
            I => n7_adj_1
        );

    \I__300\ : Odrv4
    port map (
            O => \N__2272\,
            I => n7_adj_1
        );

    \I__299\ : InMux
    port map (
            O => \N__2267\,
            I => \N__2264\
        );

    \I__298\ : LocalMux
    port map (
            O => \N__2264\,
            I => \N__2260\
        );

    \I__297\ : InMux
    port map (
            O => \N__2263\,
            I => \N__2257\
        );

    \I__296\ : Span4Mux_h
    port map (
            O => \N__2260\,
            I => \N__2254\
        );

    \I__295\ : LocalMux
    port map (
            O => \N__2257\,
            I => \ctrl_ledsArea_shifter_0\
        );

    \I__294\ : Odrv4
    port map (
            O => \N__2254\,
            I => \ctrl_ledsArea_shifter_0\
        );

    \I__293\ : CascadeMux
    port map (
            O => \N__2249\,
            I => \ctrl_tap_tdoUnbufferd_N_211_cascade_\
        );

    \I__292\ : IoInMux
    port map (
            O => \N__2246\,
            I => \N__2243\
        );

    \I__291\ : LocalMux
    port map (
            O => \N__2243\,
            I => \N__2240\
        );

    \I__290\ : Odrv12
    port map (
            O => \N__2240\,
            I => \ctrl_tap_tdoUnbufferd\
        );

    \I__289\ : InMux
    port map (
            O => \N__2237\,
            I => n2078
        );

    \I__288\ : InMux
    port map (
            O => \N__2234\,
            I => n2079
        );

    \I__287\ : InMux
    port map (
            O => \N__2231\,
            I => n2080
        );

    \I__286\ : SRMux
    port map (
            O => \N__2228\,
            I => \N__2224\
        );

    \I__285\ : SRMux
    port map (
            O => \N__2227\,
            I => \N__2220\
        );

    \I__284\ : LocalMux
    port map (
            O => \N__2224\,
            I => \N__2217\
        );

    \I__283\ : SRMux
    port map (
            O => \N__2223\,
            I => \N__2214\
        );

    \I__282\ : LocalMux
    port map (
            O => \N__2220\,
            I => \N__2210\
        );

    \I__281\ : Span4Mux_v
    port map (
            O => \N__2217\,
            I => \N__2205\
        );

    \I__280\ : LocalMux
    port map (
            O => \N__2214\,
            I => \N__2205\
        );

    \I__279\ : SRMux
    port map (
            O => \N__2213\,
            I => \N__2202\
        );

    \I__278\ : Span4Mux_v
    port map (
            O => \N__2210\,
            I => \N__2195\
        );

    \I__277\ : Span4Mux_h
    port map (
            O => \N__2205\,
            I => \N__2195\
        );

    \I__276\ : LocalMux
    port map (
            O => \N__2202\,
            I => \N__2195\
        );

    \I__275\ : Span4Mux_v
    port map (
            O => \N__2195\,
            I => \N__2192\
        );

    \I__274\ : IoSpan4Mux
    port map (
            O => \N__2192\,
            I => \N__2189\
        );

    \I__273\ : Odrv4
    port map (
            O => \N__2189\,
            I => global_reset_c
        );

    \I__272\ : InMux
    port map (
            O => \N__2186\,
            I => \N__2180\
        );

    \I__271\ : InMux
    port map (
            O => \N__2185\,
            I => \N__2180\
        );

    \I__270\ : LocalMux
    port map (
            O => \N__2180\,
            I => \ctrl_idcodeArea_shifter_31\
        );

    \I__269\ : InMux
    port map (
            O => \N__2177\,
            I => \N__2171\
        );

    \I__268\ : InMux
    port map (
            O => \N__2176\,
            I => \N__2171\
        );

    \I__267\ : LocalMux
    port map (
            O => \N__2171\,
            I => \ctrl_idcodeArea_shifter_28\
        );

    \I__266\ : CascadeMux
    port map (
            O => \N__2168\,
            I => \N__2165\
        );

    \I__265\ : InMux
    port map (
            O => \N__2165\,
            I => \N__2159\
        );

    \I__264\ : InMux
    port map (
            O => \N__2164\,
            I => \N__2159\
        );

    \I__263\ : LocalMux
    port map (
            O => \N__2159\,
            I => \ctrl_idcodeArea_shifter_30\
        );

    \I__262\ : InMux
    port map (
            O => \N__2156\,
            I => \N__2150\
        );

    \I__261\ : InMux
    port map (
            O => \N__2155\,
            I => \N__2150\
        );

    \I__260\ : LocalMux
    port map (
            O => \N__2150\,
            I => \ctrl_idcodeArea_shifter_29\
        );

    \I__259\ : InMux
    port map (
            O => \N__2147\,
            I => n2069
        );

    \I__258\ : InMux
    port map (
            O => \N__2144\,
            I => n2070
        );

    \I__257\ : InMux
    port map (
            O => \N__2141\,
            I => n2071
        );

    \I__256\ : InMux
    port map (
            O => \N__2138\,
            I => n2072
        );

    \I__255\ : InMux
    port map (
            O => \N__2135\,
            I => n2073
        );

    \I__254\ : InMux
    port map (
            O => \N__2132\,
            I => \bfn_4_9_0_\
        );

    \I__253\ : InMux
    port map (
            O => \N__2129\,
            I => n2075
        );

    \I__252\ : InMux
    port map (
            O => \N__2126\,
            I => n2076
        );

    \I__251\ : InMux
    port map (
            O => \N__2123\,
            I => n2077
        );

    \I__250\ : InMux
    port map (
            O => \N__2120\,
            I => n2060
        );

    \I__249\ : InMux
    port map (
            O => \N__2117\,
            I => n2061
        );

    \I__248\ : InMux
    port map (
            O => \N__2114\,
            I => n2062
        );

    \I__247\ : InMux
    port map (
            O => \N__2111\,
            I => n2063
        );

    \I__246\ : InMux
    port map (
            O => \N__2108\,
            I => n2064
        );

    \I__245\ : InMux
    port map (
            O => \N__2105\,
            I => n2065
        );

    \I__244\ : InMux
    port map (
            O => \N__2102\,
            I => \bfn_4_8_0_\
        );

    \I__243\ : InMux
    port map (
            O => \N__2099\,
            I => n2067
        );

    \I__242\ : InMux
    port map (
            O => \N__2096\,
            I => n2068
        );

    \I__241\ : InMux
    port map (
            O => \N__2093\,
            I => \N__2090\
        );

    \I__240\ : LocalMux
    port map (
            O => \N__2090\,
            I => \N__2087\
        );

    \I__239\ : Odrv4
    port map (
            O => \N__2087\,
            I => n7
        );

    \I__238\ : CascadeMux
    port map (
            O => \N__2084\,
            I => \n7_cascade_\
        );

    \I__237\ : InMux
    port map (
            O => \N__2081\,
            I => \N__2078\
        );

    \I__236\ : LocalMux
    port map (
            O => \N__2078\,
            I => n2206
        );

    \I__235\ : CascadeMux
    port map (
            O => \N__2075\,
            I => \n7_adj_1_cascade_\
        );

    \I__234\ : InMux
    port map (
            O => \N__2072\,
            I => \bfn_4_7_0_\
        );

    \I__233\ : InMux
    port map (
            O => \N__2069\,
            I => n2059
        );

    \I__232\ : InMux
    port map (
            O => \N__2066\,
            I => \N__2060\
        );

    \I__231\ : InMux
    port map (
            O => \N__2065\,
            I => \N__2060\
        );

    \I__230\ : LocalMux
    port map (
            O => \N__2060\,
            I => \ctrl_idcodeArea_shifter_16\
        );

    \I__229\ : CascadeMux
    port map (
            O => \N__2057\,
            I => \N__2053\
        );

    \I__228\ : CascadeMux
    port map (
            O => \N__2056\,
            I => \N__2050\
        );

    \I__227\ : InMux
    port map (
            O => \N__2053\,
            I => \N__2045\
        );

    \I__226\ : InMux
    port map (
            O => \N__2050\,
            I => \N__2045\
        );

    \I__225\ : LocalMux
    port map (
            O => \N__2045\,
            I => \ctrl_idcodeArea_shifter_15\
        );

    \I__224\ : CascadeMux
    port map (
            O => \N__2042\,
            I => \N__2038\
        );

    \I__223\ : InMux
    port map (
            O => \N__2041\,
            I => \N__2033\
        );

    \I__222\ : InMux
    port map (
            O => \N__2038\,
            I => \N__2033\
        );

    \I__221\ : LocalMux
    port map (
            O => \N__2033\,
            I => \ctrl_idcodeArea_shifter_14\
        );

    \I__220\ : CascadeMux
    port map (
            O => \N__2030\,
            I => \N__2026\
        );

    \I__219\ : InMux
    port map (
            O => \N__2029\,
            I => \N__2021\
        );

    \I__218\ : InMux
    port map (
            O => \N__2026\,
            I => \N__2021\
        );

    \I__217\ : LocalMux
    port map (
            O => \N__2021\,
            I => \ctrl_idcodeArea_shifter_13\
        );

    \I__216\ : CascadeMux
    port map (
            O => \N__2018\,
            I => \N__2014\
        );

    \I__215\ : InMux
    port map (
            O => \N__2017\,
            I => \N__2009\
        );

    \I__214\ : InMux
    port map (
            O => \N__2014\,
            I => \N__2009\
        );

    \I__213\ : LocalMux
    port map (
            O => \N__2009\,
            I => \ctrl_idcodeArea_shifter_12\
        );

    \I__212\ : CascadeMux
    port map (
            O => \N__2006\,
            I => \N__2003\
        );

    \I__211\ : InMux
    port map (
            O => \N__2003\,
            I => \N__1999\
        );

    \I__210\ : InMux
    port map (
            O => \N__2002\,
            I => \N__1996\
        );

    \I__209\ : LocalMux
    port map (
            O => \N__1999\,
            I => \ctrl_idcodeArea_shifter_3\
        );

    \I__208\ : LocalMux
    port map (
            O => \N__1996\,
            I => \ctrl_idcodeArea_shifter_3\
        );

    \I__207\ : CascadeMux
    port map (
            O => \N__1991\,
            I => \N__1987\
        );

    \I__206\ : CascadeMux
    port map (
            O => \N__1990\,
            I => \N__1984\
        );

    \I__205\ : InMux
    port map (
            O => \N__1987\,
            I => \N__1979\
        );

    \I__204\ : InMux
    port map (
            O => \N__1984\,
            I => \N__1979\
        );

    \I__203\ : LocalMux
    port map (
            O => \N__1979\,
            I => \ctrl_idcodeArea_shifter_2\
        );

    \I__202\ : InMux
    port map (
            O => \N__1976\,
            I => \N__1970\
        );

    \I__201\ : InMux
    port map (
            O => \N__1975\,
            I => \N__1970\
        );

    \I__200\ : LocalMux
    port map (
            O => \N__1970\,
            I => \ctrl_idcodeArea_shifter_7\
        );

    \I__199\ : CascadeMux
    port map (
            O => \N__1967\,
            I => \N__1963\
        );

    \I__198\ : InMux
    port map (
            O => \N__1966\,
            I => \N__1958\
        );

    \I__197\ : InMux
    port map (
            O => \N__1963\,
            I => \N__1958\
        );

    \I__196\ : LocalMux
    port map (
            O => \N__1958\,
            I => \ctrl_idcodeArea_shifter_10\
        );

    \I__195\ : InMux
    port map (
            O => \N__1955\,
            I => \N__1949\
        );

    \I__194\ : InMux
    port map (
            O => \N__1954\,
            I => \N__1949\
        );

    \I__193\ : LocalMux
    port map (
            O => \N__1949\,
            I => \ctrl_idcodeArea_shifter_9\
        );

    \I__192\ : InMux
    port map (
            O => \N__1946\,
            I => \N__1940\
        );

    \I__191\ : InMux
    port map (
            O => \N__1945\,
            I => \N__1940\
        );

    \I__190\ : LocalMux
    port map (
            O => \N__1940\,
            I => \ctrl_idcodeArea_shifter_8\
        );

    \I__189\ : InMux
    port map (
            O => \N__1937\,
            I => \N__1931\
        );

    \I__188\ : InMux
    port map (
            O => \N__1936\,
            I => \N__1931\
        );

    \I__187\ : LocalMux
    port map (
            O => \N__1931\,
            I => \ctrl_idcodeArea_shifter_4\
        );

    \I__186\ : CascadeMux
    port map (
            O => \N__1928\,
            I => \N__1925\
        );

    \I__185\ : InMux
    port map (
            O => \N__1925\,
            I => \N__1919\
        );

    \I__184\ : InMux
    port map (
            O => \N__1924\,
            I => \N__1919\
        );

    \I__183\ : LocalMux
    port map (
            O => \N__1919\,
            I => \ctrl_idcodeArea_shifter_6\
        );

    \I__182\ : InMux
    port map (
            O => \N__1916\,
            I => \N__1910\
        );

    \I__181\ : InMux
    port map (
            O => \N__1915\,
            I => \N__1910\
        );

    \I__180\ : LocalMux
    port map (
            O => \N__1910\,
            I => \ctrl_idcodeArea_shifter_5\
        );

    \I__179\ : CascadeMux
    port map (
            O => \N__1907\,
            I => \N__1903\
        );

    \I__178\ : InMux
    port map (
            O => \N__1906\,
            I => \N__1900\
        );

    \I__177\ : InMux
    port map (
            O => \N__1903\,
            I => \N__1897\
        );

    \I__176\ : LocalMux
    port map (
            O => \N__1900\,
            I => \ctrl_idcodeArea_shifter_11\
        );

    \I__175\ : LocalMux
    port map (
            O => \N__1897\,
            I => \ctrl_idcodeArea_shifter_11\
        );

    \I__174\ : IoInMux
    port map (
            O => \N__1892\,
            I => \N__1889\
        );

    \I__173\ : LocalMux
    port map (
            O => \N__1889\,
            I => \N__1886\
        );

    \I__172\ : IoSpan4Mux
    port map (
            O => \N__1886\,
            I => \N__1883\
        );

    \I__171\ : IoSpan4Mux
    port map (
            O => \N__1883\,
            I => \N__1880\
        );

    \I__170\ : Span4Mux_s3_h
    port map (
            O => \N__1880\,
            I => \N__1876\
        );

    \I__169\ : CascadeMux
    port map (
            O => \N__1879\,
            I => \N__1873\
        );

    \I__168\ : Sp12to4
    port map (
            O => \N__1876\,
            I => \N__1869\
        );

    \I__167\ : InMux
    port map (
            O => \N__1873\,
            I => \N__1866\
        );

    \I__166\ : InMux
    port map (
            O => \N__1872\,
            I => \N__1863\
        );

    \I__165\ : Odrv12
    port map (
            O => \N__1869\,
            I => io_leds_c_0
        );

    \I__164\ : LocalMux
    port map (
            O => \N__1866\,
            I => io_leds_c_0
        );

    \I__163\ : LocalMux
    port map (
            O => \N__1863\,
            I => io_leds_c_0
        );

    \I__162\ : IoInMux
    port map (
            O => \N__1856\,
            I => \N__1853\
        );

    \I__161\ : LocalMux
    port map (
            O => \N__1853\,
            I => \N__1850\
        );

    \I__160\ : Span4Mux_s3_h
    port map (
            O => \N__1850\,
            I => \N__1847\
        );

    \I__159\ : Span4Mux_v
    port map (
            O => \N__1847\,
            I => \N__1844\
        );

    \I__158\ : Sp12to4
    port map (
            O => \N__1844\,
            I => \N__1841\
        );

    \I__157\ : Odrv12
    port map (
            O => \N__1841\,
            I => io_jtag_tck_pad_gb_input
        );

    \IN_MUX_bfv_4_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_7_0_\
        );

    \IN_MUX_bfv_4_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n2066,
            carryinitout => \bfn_4_8_0_\
        );

    \IN_MUX_bfv_4_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n2074,
            carryinitout => \bfn_4_9_0_\
        );

    \io_jtag_tck_pad_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__1856\,
            GLOBALBUFFEROUTPUT => io_jtag_tck_c
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \ctrl_ledsArea_store_i0_i1_LC_2_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__1872\,
            in1 => \N__4415\,
            in2 => \_gnd_net_\,
            in3 => \N__2263\,
            lcout => io_leds_c_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4306\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_ledsArea_shifter_i0_i0_LC_2_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__4739\,
            in1 => \N__2093\,
            in2 => \N__1879\,
            in3 => \N__4571\,
            lcout => \ctrl_ledsArea_shifter_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4305\,
            ce => \N__4498\,
            sr => \_gnd_net_\
        );

    \ctrl_idcodeArea_shifter_i6_LC_4_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010001000"
        )
    port map (
            in0 => \N__1975\,
            in1 => \N__3278\,
            in2 => \N__1928\,
            in3 => \N__3423\,
            lcout => \ctrl_idcodeArea_shifter_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4316\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_idcodeArea_shifter_i4_LC_4_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101000010000000"
        )
    port map (
            in0 => \N__3421\,
            in1 => \N__1937\,
            in2 => \N__3295\,
            in3 => \N__1915\,
            lcout => \ctrl_idcodeArea_shifter_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4316\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_idcodeArea_shifter_i10_LC_4_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011000000"
        )
    port map (
            in0 => \N__1966\,
            in1 => \N__3270\,
            in2 => \N__1907\,
            in3 => \N__3419\,
            lcout => \ctrl_idcodeArea_shifter_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4316\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_idcodeArea_shifter_i7_LC_4_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101000010000000"
        )
    port map (
            in0 => \N__3424\,
            in1 => \N__1976\,
            in2 => \N__3297\,
            in3 => \N__1945\,
            lcout => \ctrl_idcodeArea_shifter_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4316\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_idcodeArea_shifter_i9_LC_4_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101111110011"
        )
    port map (
            in0 => \N__1955\,
            in1 => \N__3285\,
            in2 => \N__1967\,
            in3 => \N__3426\,
            lcout => \ctrl_idcodeArea_shifter_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4316\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_idcodeArea_shifter_i8_LC_4_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101111110001111"
        )
    port map (
            in0 => \N__3425\,
            in1 => \N__1946\,
            in2 => \N__3298\,
            in3 => \N__1954\,
            lcout => \ctrl_idcodeArea_shifter_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4316\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_idcodeArea_shifter_i3_LC_4_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010001000"
        )
    port map (
            in0 => \N__1936\,
            in1 => \N__3271\,
            in2 => \N__2006\,
            in3 => \N__3420\,
            lcout => \ctrl_idcodeArea_shifter_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4316\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_idcodeArea_shifter_i5_LC_4_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101111110001111"
        )
    port map (
            in0 => \N__3422\,
            in1 => \N__1916\,
            in2 => \N__3296\,
            in3 => \N__1924\,
            lcout => \ctrl_idcodeArea_shifter_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4316\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_idcodeArea_shifter_i11_LC_4_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011000000"
        )
    port map (
            in0 => \N__1906\,
            in1 => \N__3237\,
            in2 => \N__2018\,
            in3 => \N__3401\,
            lcout => \ctrl_idcodeArea_shifter_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4312\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_idcodeArea_shifter_i1_LC_4_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100000000000"
        )
    port map (
            in0 => \N__3407\,
            in1 => \N__2318\,
            in2 => \N__1990\,
            in3 => \N__3243\,
            lcout => \ctrl_idcodeArea_shifter_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4312\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_idcodeArea_shifter_i13_LC_4_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011000000"
        )
    port map (
            in0 => \N__2029\,
            in1 => \N__3239\,
            in2 => \N__2042\,
            in3 => \N__3403\,
            lcout => \ctrl_idcodeArea_shifter_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4312\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_idcodeArea_shifter_i15_LC_4_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010000000000"
        )
    port map (
            in0 => \N__3405\,
            in1 => \N__2065\,
            in2 => \N__2057\,
            in3 => \N__3242\,
            lcout => \ctrl_idcodeArea_shifter_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4312\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_idcodeArea_shifter_i16_LC_4_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101111110011"
        )
    port map (
            in0 => \N__2066\,
            in1 => \N__3240\,
            in2 => \N__2336\,
            in3 => \N__3406\,
            lcout => \ctrl_idcodeArea_shifter_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4312\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_idcodeArea_shifter_i14_LC_4_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011111111"
        )
    port map (
            in0 => \N__3404\,
            in1 => \N__2041\,
            in2 => \N__2056\,
            in3 => \N__3241\,
            lcout => \ctrl_idcodeArea_shifter_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4312\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_idcodeArea_shifter_i12_LC_4_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011000000"
        )
    port map (
            in0 => \N__2017\,
            in1 => \N__3238\,
            in2 => \N__2030\,
            in3 => \N__3402\,
            lcout => \ctrl_idcodeArea_shifter_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4312\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_idcodeArea_shifter_i2_LC_4_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010000000000"
        )
    port map (
            in0 => \N__3408\,
            in1 => \N__2002\,
            in2 => \N__1991\,
            in3 => \N__3244\,
            lcout => \ctrl_idcodeArea_shifter_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4312\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1546_2_lut_3_lut_LC_4_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011101110"
        )
    port map (
            in0 => \N__3819\,
            in1 => \N__3912\,
            in2 => \_gnd_net_\,
            in3 => \N__3721\,
            lcout => n2248,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1457_2_lut_LC_4_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3703\,
            in2 => \_gnd_net_\,
            in3 => \N__3818\,
            lcout => n2206,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1555_2_lut_LC_4_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4199\,
            in2 => \_gnd_net_\,
            in3 => \N__3722\,
            lcout => n2306,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_tap_instructionShift_i0_i0_LC_4_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__2389\,
            in1 => \N__2521\,
            in2 => \_gnd_net_\,
            in3 => \N__3704\,
            lcout => \ctrl_tap_instructionShift_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4309\,
            ce => \N__2566\,
            sr => \_gnd_net_\
        );

    \ctrl_tap_instructionShift_i0_i1_LC_4_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__2443\,
            in1 => \N__2377\,
            in2 => \_gnd_net_\,
            in3 => \N__3723\,
            lcout => \ctrl_tap_instructionShift_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4309\,
            ce => \N__2566\,
            sr => \_gnd_net_\
        );

    \ctrl_tap_instructionShift_i0_i2_LC_4_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__2491\,
            in1 => \N__2431\,
            in2 => \_gnd_net_\,
            in3 => \N__3705\,
            lcout => \ctrl_tap_instructionShift_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4309\,
            ce => \N__2566\,
            sr => \_gnd_net_\
        );

    \ctrl_tap_instructionShift_i0_i3_LC_4_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__3522\,
            in1 => \N__2480\,
            in2 => \_gnd_net_\,
            in3 => \N__3724\,
            lcout => \ctrl_tap_instructionShift_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4309\,
            ce => \N__2566\,
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_4_lut_adj_2_LC_4_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111111111"
        )
    port map (
            in0 => \N__3715\,
            in1 => \N__4034\,
            in2 => \N__4160\,
            in3 => \N__3837\,
            lcout => n7,
            ltout => \n7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_ledsArea_shifter_i0_i7_LC_4_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010101010"
        )
    port map (
            in0 => \N__3524\,
            in1 => \N__2796\,
            in2 => \N__2084\,
            in3 => \N__4570\,
            lcout => \ctrl_ledsArea_shifter_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4307\,
            ce => \N__4497\,
            sr => \_gnd_net_\
        );

    \i1_2_lut_4_lut_LC_4_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__3836\,
            in1 => \N__4156\,
            in2 => \N__2285\,
            in3 => \N__4035\,
            lcout => n1275,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_4_lut_LC_4_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111111111111"
        )
    port map (
            in0 => \N__2520\,
            in1 => \N__2474\,
            in2 => \N__2378\,
            in3 => \N__2430\,
            lcout => n7_adj_1,
            ltout => \n7_adj_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i4_4_lut_LC_4_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__4033\,
            in1 => \N__2081\,
            in2 => \N__2075\,
            in3 => \N__4155\,
            lcout => n2110,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \myClockArea_timeout_counter_value_317__i0_LC_4_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__3108\,
            in1 => \N__2738\,
            in2 => \_gnd_net_\,
            in3 => \N__2072\,
            lcout => \myClockArea_timeout_counter_value_0\,
            ltout => OPEN,
            carryin => \bfn_4_7_0_\,
            carryout => n2059,
            clk => \N__2846\,
            ce => 'H',
            sr => \N__2227\
        );

    \myClockArea_timeout_counter_value_317__i1_LC_4_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__3095\,
            in1 => \N__2765\,
            in2 => \_gnd_net_\,
            in3 => \N__2069\,
            lcout => \myClockArea_timeout_counter_value_1\,
            ltout => OPEN,
            carryin => n2059,
            carryout => n2060,
            clk => \N__2846\,
            ce => 'H',
            sr => \N__2227\
        );

    \myClockArea_timeout_counter_value_317__i2_LC_4_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__3109\,
            in1 => \N__2630\,
            in2 => \_gnd_net_\,
            in3 => \N__2120\,
            lcout => \myClockArea_timeout_counter_value_2\,
            ltout => OPEN,
            carryin => n2060,
            carryout => n2061,
            clk => \N__2846\,
            ce => 'H',
            sr => \N__2227\
        );

    \myClockArea_timeout_counter_value_317__i3_LC_4_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__3096\,
            in1 => \N__2777\,
            in2 => \_gnd_net_\,
            in3 => \N__2117\,
            lcout => \myClockArea_timeout_counter_value_3\,
            ltout => OPEN,
            carryin => n2061,
            carryout => n2062,
            clk => \N__2846\,
            ce => 'H',
            sr => \N__2227\
        );

    \myClockArea_timeout_counter_value_317__i4_LC_4_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__3110\,
            in1 => \N__2720\,
            in2 => \_gnd_net_\,
            in3 => \N__2114\,
            lcout => \myClockArea_timeout_counter_value_4\,
            ltout => OPEN,
            carryin => n2062,
            carryout => n2063,
            clk => \N__2846\,
            ce => 'H',
            sr => \N__2227\
        );

    \myClockArea_timeout_counter_value_317__i5_LC_4_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__3097\,
            in1 => \N__2752\,
            in2 => \_gnd_net_\,
            in3 => \N__2111\,
            lcout => \myClockArea_timeout_counter_value_5\,
            ltout => OPEN,
            carryin => n2063,
            carryout => n2064,
            clk => \N__2846\,
            ce => 'H',
            sr => \N__2227\
        );

    \myClockArea_timeout_counter_value_317__i6_LC_4_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__3111\,
            in1 => \N__2708\,
            in2 => \_gnd_net_\,
            in3 => \N__2108\,
            lcout => \myClockArea_timeout_counter_value_6\,
            ltout => OPEN,
            carryin => n2064,
            carryout => n2065,
            clk => \N__2846\,
            ce => 'H',
            sr => \N__2227\
        );

    \myClockArea_timeout_counter_value_317__i7_LC_4_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__3098\,
            in1 => \N__3029\,
            in2 => \_gnd_net_\,
            in3 => \N__2105\,
            lcout => \myClockArea_timeout_counter_value_7\,
            ltout => OPEN,
            carryin => n2065,
            carryout => n2066,
            clk => \N__2846\,
            ce => 'H',
            sr => \N__2227\
        );

    \myClockArea_timeout_counter_value_317__i8_LC_4_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__3119\,
            in1 => \N__2657\,
            in2 => \_gnd_net_\,
            in3 => \N__2102\,
            lcout => \myClockArea_timeout_counter_value_8\,
            ltout => OPEN,
            carryin => \bfn_4_8_0_\,
            carryout => n2067,
            clk => \N__2845\,
            ce => 'H',
            sr => \N__2228\
        );

    \myClockArea_timeout_counter_value_317__i9_LC_4_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__3091\,
            in1 => \N__2942\,
            in2 => \_gnd_net_\,
            in3 => \N__2099\,
            lcout => \myClockArea_timeout_counter_value_9\,
            ltout => OPEN,
            carryin => n2067,
            carryout => n2068,
            clk => \N__2845\,
            ce => 'H',
            sr => \N__2228\
        );

    \myClockArea_timeout_counter_value_317__i10_LC_4_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__3116\,
            in1 => \N__2644\,
            in2 => \_gnd_net_\,
            in3 => \N__2096\,
            lcout => \myClockArea_timeout_counter_value_10\,
            ltout => OPEN,
            carryin => n2068,
            carryout => n2069,
            clk => \N__2845\,
            ce => 'H',
            sr => \N__2228\
        );

    \myClockArea_timeout_counter_value_317__i11_LC_4_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__3088\,
            in1 => \N__2960\,
            in2 => \_gnd_net_\,
            in3 => \N__2147\,
            lcout => \myClockArea_timeout_counter_value_11\,
            ltout => OPEN,
            carryin => n2069,
            carryout => n2070,
            clk => \N__2845\,
            ce => 'H',
            sr => \N__2228\
        );

    \myClockArea_timeout_counter_value_317__i12_LC_4_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__3117\,
            in1 => \N__2917\,
            in2 => \_gnd_net_\,
            in3 => \N__2144\,
            lcout => \myClockArea_timeout_counter_value_12\,
            ltout => OPEN,
            carryin => n2070,
            carryout => n2071,
            clk => \N__2845\,
            ce => 'H',
            sr => \N__2228\
        );

    \myClockArea_timeout_counter_value_317__i13_LC_4_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__3089\,
            in1 => \N__2603\,
            in2 => \_gnd_net_\,
            in3 => \N__2141\,
            lcout => \myClockArea_timeout_counter_value_13\,
            ltout => OPEN,
            carryin => n2071,
            carryout => n2072,
            clk => \N__2845\,
            ce => 'H',
            sr => \N__2228\
        );

    \myClockArea_timeout_counter_value_317__i14_LC_4_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__3118\,
            in1 => \N__2903\,
            in2 => \_gnd_net_\,
            in3 => \N__2138\,
            lcout => \myClockArea_timeout_counter_value_14\,
            ltout => OPEN,
            carryin => n2072,
            carryout => n2073,
            clk => \N__2845\,
            ce => 'H',
            sr => \N__2228\
        );

    \myClockArea_timeout_counter_value_317__i15_LC_4_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__3090\,
            in1 => \N__2987\,
            in2 => \_gnd_net_\,
            in3 => \N__2135\,
            lcout => \myClockArea_timeout_counter_value_15\,
            ltout => OPEN,
            carryin => n2073,
            carryout => n2074,
            clk => \N__2845\,
            ce => 'H',
            sr => \N__2228\
        );

    \myClockArea_timeout_counter_value_317__i16_LC_4_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__3112\,
            in1 => \N__2681\,
            in2 => \_gnd_net_\,
            in3 => \N__2132\,
            lcout => \myClockArea_timeout_counter_value_16\,
            ltout => OPEN,
            carryin => \bfn_4_9_0_\,
            carryout => n2075,
            clk => \N__2847\,
            ce => 'H',
            sr => \N__2223\
        );

    \myClockArea_timeout_counter_value_317__i17_LC_4_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__3092\,
            in1 => \N__2669\,
            in2 => \_gnd_net_\,
            in3 => \N__2129\,
            lcout => \myClockArea_timeout_counter_value_17\,
            ltout => OPEN,
            carryin => n2075,
            carryout => n2076,
            clk => \N__2847\,
            ce => 'H',
            sr => \N__2223\
        );

    \myClockArea_timeout_counter_value_317__i18_LC_4_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__3113\,
            in1 => \N__2930\,
            in2 => \_gnd_net_\,
            in3 => \N__2126\,
            lcout => \myClockArea_timeout_counter_value_18\,
            ltout => OPEN,
            carryin => n2076,
            carryout => n2077,
            clk => \N__2847\,
            ce => 'H',
            sr => \N__2223\
        );

    \myClockArea_timeout_counter_value_317__i19_LC_4_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__3093\,
            in1 => \N__2999\,
            in2 => \_gnd_net_\,
            in3 => \N__2123\,
            lcout => \myClockArea_timeout_counter_value_19\,
            ltout => OPEN,
            carryin => n2077,
            carryout => n2078,
            clk => \N__2847\,
            ce => 'H',
            sr => \N__2223\
        );

    \myClockArea_timeout_counter_value_317__i20_LC_4_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__3114\,
            in1 => \N__2974\,
            in2 => \_gnd_net_\,
            in3 => \N__2237\,
            lcout => \myClockArea_timeout_counter_value_20\,
            ltout => OPEN,
            carryin => n2078,
            carryout => n2079,
            clk => \N__2847\,
            ce => 'H',
            sr => \N__2223\
        );

    \myClockArea_timeout_counter_value_317__i21_LC_4_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__3094\,
            in1 => \N__3017\,
            in2 => \_gnd_net_\,
            in3 => \N__2234\,
            lcout => \myClockArea_timeout_counter_value_21\,
            ltout => OPEN,
            carryin => n2079,
            carryout => n2080,
            clk => \N__2847\,
            ce => 'H',
            sr => \N__2223\
        );

    \myClockArea_timeout_counter_value_317__i22_LC_4_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__3115\,
            in1 => \N__2695\,
            in2 => \_gnd_net_\,
            in3 => \N__2231\,
            lcout => \myClockArea_timeout_counter_value_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2847\,
            ce => 'H',
            sr => \N__2223\
        );

    \myClockArea_timeout_state_90_LC_4_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__2588\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2883\,
            lcout => \myClockArea_timeout_state\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2848\,
            ce => 'H',
            sr => \N__2213\
        );

    \ctrl_idcodeArea_shifter_i28_LC_5_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101000010000000"
        )
    port map (
            in0 => \N__3415\,
            in1 => \N__2177\,
            in2 => \N__3292\,
            in3 => \N__2155\,
            lcout => \ctrl_idcodeArea_shifter_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4319\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_idcodeArea_shifter_i30_LC_5_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010001000"
        )
    port map (
            in0 => \N__2185\,
            in1 => \N__3266\,
            in2 => \N__2168\,
            in3 => \N__3417\,
            lcout => \ctrl_idcodeArea_shifter_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4319\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_idcodeArea_shifter_i31_LC_5_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111101001111"
        )
    port map (
            in0 => \N__3418\,
            in1 => \N__3512\,
            in2 => \N__3294\,
            in3 => \N__2186\,
            lcout => \ctrl_idcodeArea_shifter_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4319\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_idcodeArea_shifter_i27_LC_5_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010001000"
        )
    port map (
            in0 => \N__2176\,
            in1 => \N__3259\,
            in2 => \N__3554\,
            in3 => \N__3414\,
            lcout => \ctrl_idcodeArea_shifter_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4319\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_idcodeArea_shifter_i29_LC_5_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101000010000000"
        )
    port map (
            in0 => \N__3416\,
            in1 => \N__2156\,
            in2 => \N__3293\,
            in3 => \N__2164\,
            lcout => \ctrl_idcodeArea_shifter_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4319\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_idcodeArea_shifter_i17_LC_5_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100000000000"
        )
    port map (
            in0 => \N__3400\,
            in1 => \N__2332\,
            in2 => \N__3446\,
            in3 => \N__3208\,
            lcout => \ctrl_idcodeArea_shifter_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4317\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_3_lut_4_lut_adj_5_LC_5_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111111111"
        )
    port map (
            in0 => \N__2428\,
            in1 => \N__2372\,
            in2 => \N__2479\,
            in3 => \N__2518\,
            lcout => n2085,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_idcodeArea_shifter_i0_LC_5_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110011111111"
        )
    port map (
            in0 => \N__2303\,
            in1 => \N__2317\,
            in2 => \N__3431\,
            in3 => \N__3207\,
            lcout => \ctrl_idcodeArea_shifter_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4317\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_ledsArea_store_i0_i6_LC_5_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__4664\,
            in1 => \N__4677\,
            in2 => \_gnd_net_\,
            in3 => \N__4418\,
            lcout => io_leds_c_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4317\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_tap_instruction_3__I_0_i6_2_lut_LC_5_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2429\,
            in2 => \_gnd_net_\,
            in3 => \N__2470\,
            lcout => OPEN,
            ltout => \n6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \equal_316_i15_4_lut_LC_5_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__2371\,
            in1 => \N__2519\,
            in2 => \N__2306\,
            in3 => \N__4551\,
            lcout => n15,
            ltout => \n15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i397_4_lut_LC_5_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001010"
        )
    port map (
            in0 => \N__2302\,
            in1 => \N__2294\,
            in2 => \N__2288\,
            in3 => \N__3560\,
            lcout => OPEN,
            ltout => \ctrl_tap_tdoUnbufferd_N_211_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i400_4_lut_LC_5_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__2284\,
            in1 => \N__2267\,
            in2 => \N__2249\,
            in3 => \N__4552\,
            lcout => \ctrl_tap_tdoUnbufferd\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_3_lut_4_lut_adj_3_LC_5_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__3838\,
            in1 => \N__3711\,
            in2 => \N__4154\,
            in3 => \N__4039\,
            lcout => n1489,
            ltout => \n1489_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_4_lut_LC_5_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111100001111"
        )
    port map (
            in0 => \N__4040\,
            in1 => \N__3596\,
            in2 => \N__2528\,
            in3 => \N__4141\,
            lcout => n1269,
            ltout => \n1269_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_tap_instruction_i0_LC_5_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110000001100"
        )
    port map (
            in0 => \N__3206\,
            in1 => \N__2522\,
            in2 => \N__2525\,
            in3 => \N__3589\,
            lcout => ctrl_tap_instruction_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4313\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i917_4_lut_4_lut_LC_5_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000010"
        )
    port map (
            in0 => \N__4038\,
            in1 => \N__4140\,
            in2 => \N__3732\,
            in3 => \N__3839\,
            lcout => n1022,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_tap_instruction_i3_LC_5_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001010000000"
        )
    port map (
            in0 => \N__3205\,
            in1 => \N__2405\,
            in2 => \N__2495\,
            in3 => \N__2475\,
            lcout => ctrl_tap_instruction_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4313\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_tap_instruction_i2_LC_5_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110110011"
        )
    port map (
            in0 => \N__2404\,
            in1 => \N__3204\,
            in2 => \N__2447\,
            in3 => \N__2432\,
            lcout => ctrl_tap_instruction_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4313\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_tap_instruction_i1_LC_5_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001010000000"
        )
    port map (
            in0 => \N__3203\,
            in1 => \N__2403\,
            in2 => \N__2393\,
            in3 => \N__2376\,
            lcout => ctrl_tap_instruction_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4313\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_tap_fsm_state_i1_LC_5_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100000001000"
        )
    port map (
            in0 => \N__4204\,
            in1 => \N__2345\,
            in2 => \N__4235\,
            in3 => \N__3608\,
            lcout => ctrl_tap_fsm_state_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4313\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_1_LC_5_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__3821\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4120\,
            lcout => OPEN,
            ltout => \n118_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1539_2_lut_3_lut_4_lut_LC_5_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111111111"
        )
    port map (
            in0 => \N__3707\,
            in1 => \N__3952\,
            in2 => \N__2339\,
            in3 => \N__4023\,
            lcout => n2273,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1531_3_lut_4_lut_LC_5_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011101100111"
        )
    port map (
            in0 => \N__3822\,
            in1 => \N__3951\,
            in2 => \N__4042\,
            in3 => \N__4121\,
            lcout => OPEN,
            ltout => \n2282_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n2323_bdd_4_lut_LC_5_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010111000"
        )
    port map (
            in0 => \N__3746\,
            in1 => \N__2540\,
            in2 => \N__2579\,
            in3 => \N__4202\,
            lcout => OPEN,
            ltout => \n2326_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_tap_fsm_state_i0_LC_5_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000111110101"
        )
    port map (
            in0 => \N__4226\,
            in1 => \N__3950\,
            in2 => \N__2576\,
            in3 => \N__2573\,
            lcout => ctrl_tap_fsm_state_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4310\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1482_4_lut_LC_5_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110111000"
        )
    port map (
            in0 => \N__2534\,
            in1 => \N__4201\,
            in2 => \N__2567\,
            in3 => \N__4259\,
            lcout => OPEN,
            ltout => \n2231_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_tap_fsm_state_i2_LC_5_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010010100000"
        )
    port map (
            in0 => \N__4227\,
            in1 => \N__4203\,
            in2 => \N__2552\,
            in3 => \N__2549\,
            lcout => ctrl_tap_fsm_state_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4310\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n2317_bdd_4_lut_4_lut_LC_5_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110011100000"
        )
    port map (
            in0 => \N__3706\,
            in1 => \N__4022\,
            in2 => \N__4143\,
            in3 => \N__3820\,
            lcout => n1119,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1535_2_lut_3_lut_LC_5_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__4123\,
            in1 => \N__3943\,
            in2 => \_gnd_net_\,
            in3 => \N__3848\,
            lcout => OPEN,
            ltout => \n2263_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_tap_fsm_state_0__bdd_4_lut_4_lut_LC_5_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110011011000100"
        )
    port map (
            in0 => \N__4198\,
            in1 => \N__3719\,
            in2 => \N__2543\,
            in3 => \N__2726\,
            lcout => n2323,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1557_4_lut_4_lut_LC_5_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001110100010101"
        )
    port map (
            in0 => \N__4124\,
            in1 => \N__3944\,
            in2 => \N__3733\,
            in3 => \N__3849\,
            lcout => n2272,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_ledsArea_store_i0_i8_LC_5_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__4393\,
            in1 => \_gnd_net_\,
            in2 => \N__2800\,
            in3 => \N__4642\,
            lcout => io_leds_c_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4308\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1041_4_lut_4_lut_LC_5_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111101011110"
        )
    port map (
            in0 => \N__4036\,
            in1 => \N__3720\,
            in2 => \N__4144\,
            in3 => \N__3850\,
            lcout => n1117,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1473_4_lut_LC_5_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__2776\,
            in1 => \N__2764\,
            in2 => \N__2753\,
            in3 => \N__2737\,
            lcout => n2222,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1558_2_lut_LC_5_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__3945\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4122\,
            lcout => n2309,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1467_4_lut_LC_5_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__2719\,
            in1 => \N__2707\,
            in2 => \N__2696\,
            in3 => \N__2680\,
            lcout => n2216,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1469_4_lut_LC_5_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__2668\,
            in1 => \N__2656\,
            in2 => \N__2645\,
            in3 => \N__2629\,
            lcout => OPEN,
            ltout => \n2218_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1479_4_lut_LC_5_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__2618\,
            in1 => \N__2948\,
            in2 => \N__2612\,
            in3 => \N__2609\,
            lcout => OPEN,
            ltout => \n2228_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i7_4_lut_LC_5_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__2602\,
            in1 => \N__3005\,
            in2 => \N__2591\,
            in3 => \N__2891\,
            lcout => n2185,
            ltout => \n2185_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1116_2_lut_LC_5_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001010000"
        )
    port map (
            in0 => \N__2885\,
            in1 => \_gnd_net_\,
            in2 => \N__3122\,
            in3 => \_gnd_net_\,
            lcout => n1848,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i3_2_lut_LC_5_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3028\,
            in2 => \_gnd_net_\,
            in3 => \N__3016\,
            lcout => n11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1471_4_lut_LC_5_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__2998\,
            in1 => \N__2986\,
            in2 => \N__2975\,
            in3 => \N__2959\,
            lcout => n2220,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i5_4_lut_LC_5_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__2941\,
            in1 => \N__2929\,
            in2 => \N__2918\,
            in3 => \N__2902\,
            lcout => n13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_ledsArea_store_i0_i7_LC_5_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__4414\,
            in1 => \N__4582\,
            in2 => \_gnd_net_\,
            in3 => \N__4520\,
            lcout => io_leds_c_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4304\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \myClockArea_toggle_92_LC_5_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2860\,
            in2 => \_gnd_net_\,
            in3 => \N__2884\,
            lcout => io_leds_c_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2849\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_idcodeArea_shifter_i24_LC_6_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101111110001111"
        )
    port map (
            in0 => \N__3428\,
            in1 => \N__2818\,
            in2 => \N__3299\,
            in3 => \N__2827\,
            lcout => \ctrl_idcodeArea_shifter_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4321\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_idcodeArea_shifter_i25_LC_6_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101111110011"
        )
    port map (
            in0 => \N__2828\,
            in1 => \N__3290\,
            in2 => \N__3538\,
            in3 => \N__3429\,
            lcout => \ctrl_idcodeArea_shifter_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4321\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_idcodeArea_shifter_i23_LC_6_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011000000"
        )
    port map (
            in0 => \N__3484\,
            in1 => \N__3286\,
            in2 => \N__2819\,
            in3 => \N__3427\,
            lcout => \ctrl_idcodeArea_shifter_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4321\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_idcodeArea_shifter_i26_LC_6_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001110111011"
        )
    port map (
            in0 => \N__3550\,
            in1 => \N__3291\,
            in2 => \N__3539\,
            in3 => \N__3430\,
            lcout => \ctrl_idcodeArea_shifter_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4321\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_tap_bypass_83_LC_6_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3523\,
            lcout => ctrl_tap_bypass,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4320\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_idcodeArea_shifter_i20_LC_6_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010000000000"
        )
    port map (
            in0 => \N__3411\,
            in1 => \N__3454\,
            in2 => \N__3314\,
            in3 => \N__3248\,
            lcout => \ctrl_idcodeArea_shifter_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4320\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_idcodeArea_shifter_i22_LC_6_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101111110011"
        )
    port map (
            in0 => \N__3469\,
            in1 => \N__3246\,
            in2 => \N__3485\,
            in3 => \N__3413\,
            lcout => \ctrl_idcodeArea_shifter_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4320\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_idcodeArea_shifter_i21_LC_6_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011111111"
        )
    port map (
            in0 => \N__3412\,
            in1 => \N__3455\,
            in2 => \N__3470\,
            in3 => \N__3249\,
            lcout => \ctrl_idcodeArea_shifter_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4320\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1017_3_lut_4_lut_LC_6_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101001101010"
        )
    port map (
            in0 => \N__4152\,
            in1 => \N__3731\,
            in2 => \N__3949\,
            in3 => \N__3840\,
            lcout => n929,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_idcodeArea_shifter_i18_LC_6_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101111110011"
        )
    port map (
            in0 => \N__3445\,
            in1 => \N__3245\,
            in2 => \N__3134\,
            in3 => \N__3409\,
            lcout => \ctrl_idcodeArea_shifter_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4320\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_idcodeArea_shifter_i19_LC_6_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100000000000"
        )
    port map (
            in0 => \N__3410\,
            in1 => \N__3133\,
            in2 => \N__3313\,
            in3 => \N__3247\,
            lcout => \ctrl_idcodeArea_shifter_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4320\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_LC_6_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4110\,
            in2 => \_gnd_net_\,
            in3 => \N__4017\,
            lcout => n4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_adj_4_LC_6_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111010"
        )
    port map (
            in0 => \N__4021\,
            in1 => \_gnd_net_\,
            in2 => \N__3955\,
            in3 => \N__4153\,
            lcout => OPEN,
            ltout => \n17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i954_4_lut_LC_6_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000001010"
        )
    port map (
            in0 => \N__3817\,
            in1 => \N__4258\,
            in2 => \N__3614\,
            in3 => \N__3698\,
            lcout => OPEN,
            ltout => \n1687_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1485_3_lut_LC_6_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3602\,
            in2 => \N__3611\,
            in3 => \N__4200\,
            lcout => n2234,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i13_4_lut_LC_6_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__3816\,
            in1 => \N__3939\,
            in2 => \N__3730\,
            in3 => \N__4112\,
            lcout => n8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_3_lut_4_lut_LC_6_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__4111\,
            in1 => \N__3815\,
            in2 => \N__4041\,
            in3 => \N__3699\,
            lcout => n7_adj_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1449_2_lut_LC_6_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__3814\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3697\,
            lcout => n2198,
            ltout => \n2198_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1182_4_lut_LC_6_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101011001100"
        )
    port map (
            in0 => \N__3590\,
            in1 => \N__3575\,
            in2 => \N__3569\,
            in3 => \N__3566\,
            lcout => \ctrl_tap_tdoUnbufferd_N_213\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_4_lut_adj_6_LC_6_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__3841\,
            in1 => \N__3725\,
            in2 => \N__4043\,
            in3 => \N__4115\,
            lcout => n1638,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_LC_6_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__4114\,
            in1 => \N__4028\,
            in2 => \_gnd_net_\,
            in3 => \N__3842\,
            lcout => n2186,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_ledsArea_store_i0_i4_LC_6_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__4720\,
            in1 => \N__4709\,
            in2 => \_gnd_net_\,
            in3 => \N__4401\,
            lcout => \ctrl_ledsArea_store_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4314\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_4_lut_adj_7_LC_6_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__4113\,
            in1 => \N__4027\,
            in2 => \N__3851\,
            in3 => \N__3954\,
            lcout => n1686,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_ledsArea_store_i0_i2_LC_6_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__4755\,
            in1 => \N__4738\,
            in2 => \_gnd_net_\,
            in3 => \N__4400\,
            lcout => io_leds_c_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4314\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i114_3_lut_LC_6_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010111011"
        )
    port map (
            in0 => \N__3726\,
            in1 => \N__4032\,
            in2 => \_gnd_net_\,
            in3 => \N__3843\,
            lcout => OPEN,
            ltout => \n112_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1534_3_lut_LC_6_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010100000"
        )
    port map (
            in0 => \N__3953\,
            in1 => \_gnd_net_\,
            in2 => \N__4247\,
            in3 => \N__4116\,
            lcout => OPEN,
            ltout => \n2260_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_tap_fsm_state_i3_LC_6_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101111000000"
        )
    port map (
            in0 => \N__4244\,
            in1 => \N__4231\,
            in2 => \N__4208\,
            in3 => \N__4205\,
            lcout => ctrl_tap_fsm_state_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4314\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1494_3_lut_4_lut_LC_6_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111010111011"
        )
    port map (
            in0 => \N__4142\,
            in1 => \N__4037\,
            in2 => \N__3956\,
            in3 => \N__3847\,
            lcout => n2243,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_ledsArea_shifter_i0_i4_LC_7_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010001000"
        )
    port map (
            in0 => \N__4450\,
            in1 => \N__3740\,
            in2 => \N__4663\,
            in3 => \N__3734\,
            lcout => \ctrl_ledsArea_shifter_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4318\,
            ce => \N__4502\,
            sr => \_gnd_net_\
        );

    \ctrl_ledsArea_shifter_i0_i1_LC_7_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__4429\,
            in1 => \N__4624\,
            in2 => \N__4762\,
            in3 => \N__4553\,
            lcout => \ctrl_ledsArea_shifter_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4318\,
            ce => \N__4502\,
            sr => \_gnd_net_\
        );

    \ctrl_ledsArea_shifter_i0_i2_LC_7_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__4554\,
            in1 => \N__4708\,
            in2 => \N__4351\,
            in3 => \N__4627\,
            lcout => \ctrl_ledsArea_shifter_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4318\,
            ce => \N__4502\,
            sr => \_gnd_net_\
        );

    \ctrl_ledsArea_shifter_i0_i3_LC_7_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__4472\,
            in1 => \N__4625\,
            in2 => \N__4724\,
            in3 => \N__4555\,
            lcout => \ctrl_ledsArea_shifter_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4318\,
            ce => \N__4502\,
            sr => \_gnd_net_\
        );

    \ctrl_ledsArea_shifter_i0_i5_LC_7_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__4556\,
            in1 => \N__4513\,
            in2 => \N__4696\,
            in3 => \N__4628\,
            lcout => \ctrl_ledsArea_shifter_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4318\,
            ce => \N__4502\,
            sr => \_gnd_net_\
        );

    \ctrl_ledsArea_shifter_i0_i6_LC_7_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__4643\,
            in1 => \N__4626\,
            in2 => \N__4600\,
            in3 => \N__4557\,
            lcout => \ctrl_ledsArea_shifter_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4318\,
            ce => \N__4502\,
            sr => \_gnd_net_\
        );

    \ctrl_ledsArea_store_i0_i5_LC_7_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__4449\,
            in1 => \N__4471\,
            in2 => \_gnd_net_\,
            in3 => \N__4416\,
            lcout => io_leds_c_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4315\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctrl_ledsArea_store_i0_i3_LC_7_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__4338\,
            in1 => \N__4433\,
            in2 => \_gnd_net_\,
            in3 => \N__4417\,
            lcout => io_leds_c_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4311\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
